module encrypt_4pre_mix(in, out);
    input [639:0] in;
    output [639:0] out;
    wire [63:0] total;
    assign total = 0 ^ in[63:0] ^ in[127:64] ^ in[191:128] ^ in[255:192] ^ in[319:256] ^ in[383:320] ^ in[447:384] ^ in[511:448] ^ in[575:512] ^ in[639:576];
    assign out[63:0] = in[63:0] ^ total ^ (total >> 32);
    assign out[127:64] = in[127:64] ^ total ^ (total >> 32);
    assign out[191:128] = in[191:128] ^ total ^ (total >> 32);
    assign out[255:192] = in[255:192] ^ total ^ (total >> 32);
    assign out[319:256] = in[319:256] ^ total ^ (total >> 32);
    assign out[383:320] = in[383:320] ^ total ^ (total >> 32);
    assign out[447:384] = in[447:384] ^ total ^ (total >> 32);
    assign out[511:448] = in[511:448] ^ total ^ (total >> 32);
    assign out[575:512] = in[575:512] ^ total ^ (total >> 32);
    assign out[639:576] = in[639:576] ^ total ^ (total >> 32);
endmodule

module encrypt_4sbox_small0(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h3e;
        mem[1] = 6'h0a;
        mem[2] = 6'h11;
        mem[3] = 6'h26;
        mem[4] = 6'h2e;
        mem[5] = 6'h27;
        mem[6] = 6'h16;
        mem[7] = 6'h05;
        mem[8] = 6'h2a;
        mem[9] = 6'h33;
        mem[10] = 6'h06;
        mem[11] = 6'h3f;
        mem[12] = 6'h1c;
        mem[13] = 6'h0d;
        mem[14] = 6'h08;
        mem[15] = 6'h2c;
        mem[16] = 6'h32;
        mem[17] = 6'h3d;
        mem[18] = 6'h0c;
        mem[19] = 6'h21;
        mem[20] = 6'h28;
        mem[21] = 6'h0f;
        mem[22] = 6'h12;
        mem[23] = 6'h3b;
        mem[24] = 6'h3c;
        mem[25] = 6'h1b;
        mem[26] = 6'h1d;
        mem[27] = 6'h09;
        mem[28] = 6'h31;
        mem[29] = 6'h24;
        mem[30] = 6'h15;
        mem[31] = 6'h2d;
        mem[32] = 6'h0b;
        mem[33] = 6'h34;
        mem[34] = 6'h23;
        mem[35] = 6'h22;
        mem[36] = 6'h3a;
        mem[37] = 6'h10;
        mem[38] = 6'h1f;
        mem[39] = 6'h17;
        mem[40] = 6'h0e;
        mem[41] = 6'h03;
        mem[42] = 6'h30;
        mem[43] = 6'h01;
        mem[44] = 6'h18;
        mem[45] = 6'h38;
        mem[46] = 6'h19;
        mem[47] = 6'h35;
        mem[48] = 6'h14;
        mem[49] = 6'h04;
        mem[50] = 6'h36;
        mem[51] = 6'h1a;
        mem[52] = 6'h2f;
        mem[53] = 6'h39;
        mem[54] = 6'h1e;
        mem[55] = 6'h37;
        mem[56] = 6'h13;
        mem[57] = 6'h20;
        mem[58] = 6'h29;
        mem[59] = 6'h02;
        mem[60] = 6'h25;
        mem[61] = 6'h2b;
        mem[62] = 6'h00;
        mem[63] = 6'h07;
    end
endmodule

module encrypt_4sbox_small1(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h03;
        mem[1] = 6'h2e;
        mem[2] = 6'h0c;
        mem[3] = 6'h2c;
        mem[4] = 6'h15;
        mem[5] = 6'h14;
        mem[6] = 6'h3c;
        mem[7] = 6'h1c;
        mem[8] = 6'h16;
        mem[9] = 6'h0a;
        mem[10] = 6'h24;
        mem[11] = 6'h17;
        mem[12] = 6'h1a;
        mem[13] = 6'h33;
        mem[14] = 6'h27;
        mem[15] = 6'h28;
        mem[16] = 6'h3f;
        mem[17] = 6'h18;
        mem[18] = 6'h09;
        mem[19] = 6'h07;
        mem[20] = 6'h04;
        mem[21] = 6'h13;
        mem[22] = 6'h05;
        mem[23] = 6'h3e;
        mem[24] = 6'h25;
        mem[25] = 6'h00;
        mem[26] = 6'h34;
        mem[27] = 6'h0f;
        mem[28] = 6'h26;
        mem[29] = 6'h1b;
        mem[30] = 6'h3b;
        mem[31] = 6'h0e;
        mem[32] = 6'h30;
        mem[33] = 6'h2a;
        mem[34] = 6'h36;
        mem[35] = 6'h38;
        mem[36] = 6'h37;
        mem[37] = 6'h21;
        mem[38] = 6'h20;
        mem[39] = 6'h29;
        mem[40] = 6'h06;
        mem[41] = 6'h0b;
        mem[42] = 6'h22;
        mem[43] = 6'h2b;
        mem[44] = 6'h0d;
        mem[45] = 6'h2f;
        mem[46] = 6'h11;
        mem[47] = 6'h23;
        mem[48] = 6'h1e;
        mem[49] = 6'h08;
        mem[50] = 6'h39;
        mem[51] = 6'h1d;
        mem[52] = 6'h2d;
        mem[53] = 6'h01;
        mem[54] = 6'h12;
        mem[55] = 6'h35;
        mem[56] = 6'h31;
        mem[57] = 6'h19;
        mem[58] = 6'h3d;
        mem[59] = 6'h02;
        mem[60] = 6'h10;
        mem[61] = 6'h32;
        mem[62] = 6'h3a;
        mem[63] = 6'h1f;
    end
endmodule

module encrypt_4sbox_small2(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h3d;
        mem[1] = 6'h3b;
        mem[2] = 6'h21;
        mem[3] = 6'h23;
        mem[4] = 6'h0c;
        mem[5] = 6'h29;
        mem[6] = 6'h14;
        mem[7] = 6'h05;
        mem[8] = 6'h32;
        mem[9] = 6'h38;
        mem[10] = 6'h11;
        mem[11] = 6'h24;
        mem[12] = 6'h31;
        mem[13] = 6'h0f;
        mem[14] = 6'h1e;
        mem[15] = 6'h37;
        mem[16] = 6'h2b;
        mem[17] = 6'h3f;
        mem[18] = 6'h1a;
        mem[19] = 6'h02;
        mem[20] = 6'h06;
        mem[21] = 6'h27;
        mem[22] = 6'h12;
        mem[23] = 6'h1b;
        mem[24] = 6'h1f;
        mem[25] = 6'h3a;
        mem[26] = 6'h26;
        mem[27] = 6'h25;
        mem[28] = 6'h03;
        mem[29] = 6'h17;
        mem[30] = 6'h07;
        mem[31] = 6'h18;
        mem[32] = 6'h22;
        mem[33] = 6'h39;
        mem[34] = 6'h0a;
        mem[35] = 6'h0d;
        mem[36] = 6'h2a;
        mem[37] = 6'h10;
        mem[38] = 6'h2e;
        mem[39] = 6'h13;
        mem[40] = 6'h00;
        mem[41] = 6'h20;
        mem[42] = 6'h2d;
        mem[43] = 6'h19;
        mem[44] = 6'h2f;
        mem[45] = 6'h1c;
        mem[46] = 6'h04;
        mem[47] = 6'h36;
        mem[48] = 6'h0b;
        mem[49] = 6'h16;
        mem[50] = 6'h08;
        mem[51] = 6'h0e;
        mem[52] = 6'h1d;
        mem[53] = 6'h34;
        mem[54] = 6'h01;
        mem[55] = 6'h09;
        mem[56] = 6'h3e;
        mem[57] = 6'h2c;
        mem[58] = 6'h35;
        mem[59] = 6'h15;
        mem[60] = 6'h30;
        mem[61] = 6'h3c;
        mem[62] = 6'h28;
        mem[63] = 6'h33;
    end
endmodule

module encrypt_4sbox_small3(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h37;
        mem[1] = 6'h13;
        mem[2] = 6'h28;
        mem[3] = 6'h00;
        mem[4] = 6'h1b;
        mem[5] = 6'h1d;
        mem[6] = 6'h2a;
        mem[7] = 6'h21;
        mem[8] = 6'h17;
        mem[9] = 6'h04;
        mem[10] = 6'h02;
        mem[11] = 6'h08;
        mem[12] = 6'h29;
        mem[13] = 6'h3c;
        mem[14] = 6'h20;
        mem[15] = 6'h3a;
        mem[16] = 6'h2b;
        mem[17] = 6'h3b;
        mem[18] = 6'h1f;
        mem[19] = 6'h27;
        mem[20] = 6'h31;
        mem[21] = 6'h33;
        mem[22] = 6'h03;
        mem[23] = 6'h38;
        mem[24] = 6'h3f;
        mem[25] = 6'h2c;
        mem[26] = 6'h34;
        mem[27] = 6'h2d;
        mem[28] = 6'h16;
        mem[29] = 6'h1c;
        mem[30] = 6'h05;
        mem[31] = 6'h0d;
        mem[32] = 6'h26;
        mem[33] = 6'h14;
        mem[34] = 6'h0f;
        mem[35] = 6'h1a;
        mem[36] = 6'h39;
        mem[37] = 6'h07;
        mem[38] = 6'h18;
        mem[39] = 6'h36;
        mem[40] = 6'h2e;
        mem[41] = 6'h06;
        mem[42] = 6'h3e;
        mem[43] = 6'h30;
        mem[44] = 6'h0e;
        mem[45] = 6'h12;
        mem[46] = 6'h32;
        mem[47] = 6'h1e;
        mem[48] = 6'h23;
        mem[49] = 6'h3d;
        mem[50] = 6'h19;
        mem[51] = 6'h2f;
        mem[52] = 6'h24;
        mem[53] = 6'h0c;
        mem[54] = 6'h11;
        mem[55] = 6'h22;
        mem[56] = 6'h0a;
        mem[57] = 6'h10;
        mem[58] = 6'h09;
        mem[59] = 6'h0b;
        mem[60] = 6'h25;
        mem[61] = 6'h35;
        mem[62] = 6'h01;
        mem[63] = 6'h15;
    end
endmodule

module encrypt_4sbox_small4(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h3e;
        mem[1] = 6'h32;
        mem[2] = 6'h25;
        mem[3] = 6'h3b;
        mem[4] = 6'h21;
        mem[5] = 6'h0c;
        mem[6] = 6'h16;
        mem[7] = 6'h2e;
        mem[8] = 6'h05;
        mem[9] = 6'h3c;
        mem[10] = 6'h10;
        mem[11] = 6'h03;
        mem[12] = 6'h20;
        mem[13] = 6'h1a;
        mem[14] = 6'h0f;
        mem[15] = 6'h01;
        mem[16] = 6'h29;
        mem[17] = 6'h09;
        mem[18] = 6'h00;
        mem[19] = 6'h13;
        mem[20] = 6'h22;
        mem[21] = 6'h11;
        mem[22] = 6'h34;
        mem[23] = 6'h1d;
        mem[24] = 6'h1b;
        mem[25] = 6'h08;
        mem[26] = 6'h02;
        mem[27] = 6'h24;
        mem[28] = 6'h30;
        mem[29] = 6'h2f;
        mem[30] = 6'h3a;
        mem[31] = 6'h07;
        mem[32] = 6'h04;
        mem[33] = 6'h38;
        mem[34] = 6'h14;
        mem[35] = 6'h28;
        mem[36] = 6'h3f;
        mem[37] = 6'h2d;
        mem[38] = 6'h17;
        mem[39] = 6'h1f;
        mem[40] = 6'h0b;
        mem[41] = 6'h0a;
        mem[42] = 6'h37;
        mem[43] = 6'h36;
        mem[44] = 6'h1e;
        mem[45] = 6'h31;
        mem[46] = 6'h12;
        mem[47] = 6'h26;
        mem[48] = 6'h23;
        mem[49] = 6'h18;
        mem[50] = 6'h2a;
        mem[51] = 6'h0d;
        mem[52] = 6'h19;
        mem[53] = 6'h15;
        mem[54] = 6'h06;
        mem[55] = 6'h39;
        mem[56] = 6'h35;
        mem[57] = 6'h2c;
        mem[58] = 6'h1c;
        mem[59] = 6'h27;
        mem[60] = 6'h2b;
        mem[61] = 6'h33;
        mem[62] = 6'h3d;
        mem[63] = 6'h0e;
    end
endmodule

module encrypt_4sbox_small5(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h0a;
        mem[1] = 6'h1b;
        mem[2] = 6'h08;
        mem[3] = 6'h03;
        mem[4] = 6'h26;
        mem[5] = 6'h3c;
        mem[6] = 6'h3d;
        mem[7] = 6'h06;
        mem[8] = 6'h38;
        mem[9] = 6'h37;
        mem[10] = 6'h10;
        mem[11] = 6'h0f;
        mem[12] = 6'h11;
        mem[13] = 6'h12;
        mem[14] = 6'h32;
        mem[15] = 6'h34;
        mem[16] = 6'h1f;
        mem[17] = 6'h30;
        mem[18] = 6'h3f;
        mem[19] = 6'h36;
        mem[20] = 6'h14;
        mem[21] = 6'h28;
        mem[22] = 6'h16;
        mem[23] = 6'h09;
        mem[24] = 6'h2c;
        mem[25] = 6'h18;
        mem[26] = 6'h3e;
        mem[27] = 6'h2d;
        mem[28] = 6'h31;
        mem[29] = 6'h19;
        mem[30] = 6'h24;
        mem[31] = 6'h0d;
        mem[32] = 6'h0e;
        mem[33] = 6'h07;
        mem[34] = 6'h2a;
        mem[35] = 6'h1a;
        mem[36] = 6'h29;
        mem[37] = 6'h2f;
        mem[38] = 6'h3a;
        mem[39] = 6'h22;
        mem[40] = 6'h2e;
        mem[41] = 6'h1e;
        mem[42] = 6'h39;
        mem[43] = 6'h2b;
        mem[44] = 6'h00;
        mem[45] = 6'h13;
        mem[46] = 6'h04;
        mem[47] = 6'h01;
        mem[48] = 6'h35;
        mem[49] = 6'h1d;
        mem[50] = 6'h20;
        mem[51] = 6'h27;
        mem[52] = 6'h05;
        mem[53] = 6'h21;
        mem[54] = 6'h25;
        mem[55] = 6'h1c;
        mem[56] = 6'h0c;
        mem[57] = 6'h23;
        mem[58] = 6'h17;
        mem[59] = 6'h15;
        mem[60] = 6'h02;
        mem[61] = 6'h3b;
        mem[62] = 6'h0b;
        mem[63] = 6'h33;
    end
endmodule

module encrypt_4sbox_small6(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h35;
        mem[1] = 6'h38;
        mem[2] = 6'h22;
        mem[3] = 6'h30;
        mem[4] = 6'h2a;
        mem[5] = 6'h15;
        mem[6] = 6'h0b;
        mem[7] = 6'h26;
        mem[8] = 6'h2f;
        mem[9] = 6'h23;
        mem[10] = 6'h0f;
        mem[11] = 6'h17;
        mem[12] = 6'h13;
        mem[13] = 6'h0c;
        mem[14] = 6'h33;
        mem[15] = 6'h24;
        mem[16] = 6'h2c;
        mem[17] = 6'h09;
        mem[18] = 6'h07;
        mem[19] = 6'h36;
        mem[20] = 6'h02;
        mem[21] = 6'h21;
        mem[22] = 6'h0d;
        mem[23] = 6'h3d;
        mem[24] = 6'h32;
        mem[25] = 6'h18;
        mem[26] = 6'h39;
        mem[27] = 6'h20;
        mem[28] = 6'h3f;
        mem[29] = 6'h3e;
        mem[30] = 6'h1e;
        mem[31] = 6'h16;
        mem[32] = 6'h2d;
        mem[33] = 6'h12;
        mem[34] = 6'h25;
        mem[35] = 6'h00;
        mem[36] = 6'h1b;
        mem[37] = 6'h1f;
        mem[38] = 6'h31;
        mem[39] = 6'h10;
        mem[40] = 6'h29;
        mem[41] = 6'h03;
        mem[42] = 6'h37;
        mem[43] = 6'h0e;
        mem[44] = 6'h05;
        mem[45] = 6'h0a;
        mem[46] = 6'h01;
        mem[47] = 6'h1a;
        mem[48] = 6'h06;
        mem[49] = 6'h2e;
        mem[50] = 6'h2b;
        mem[51] = 6'h1d;
        mem[52] = 6'h3b;
        mem[53] = 6'h3c;
        mem[54] = 6'h19;
        mem[55] = 6'h08;
        mem[56] = 6'h04;
        mem[57] = 6'h1c;
        mem[58] = 6'h14;
        mem[59] = 6'h28;
        mem[60] = 6'h11;
        mem[61] = 6'h34;
        mem[62] = 6'h27;
        mem[63] = 6'h3a;
    end
endmodule

module encrypt_4sbox_small7(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h32;
        mem[1] = 6'h2a;
        mem[2] = 6'h20;
        mem[3] = 6'h1a;
        mem[4] = 6'h2f;
        mem[5] = 6'h18;
        mem[6] = 6'h16;
        mem[7] = 6'h11;
        mem[8] = 6'h2d;
        mem[9] = 6'h22;
        mem[10] = 6'h29;
        mem[11] = 6'h23;
        mem[12] = 6'h37;
        mem[13] = 6'h04;
        mem[14] = 6'h2b;
        mem[15] = 6'h38;
        mem[16] = 6'h2c;
        mem[17] = 6'h1c;
        mem[18] = 6'h13;
        mem[19] = 6'h33;
        mem[20] = 6'h39;
        mem[21] = 6'h19;
        mem[22] = 6'h0c;
        mem[23] = 6'h24;
        mem[24] = 6'h1e;
        mem[25] = 6'h3d;
        mem[26] = 6'h02;
        mem[27] = 6'h26;
        mem[28] = 6'h27;
        mem[29] = 6'h1f;
        mem[30] = 6'h14;
        mem[31] = 6'h31;
        mem[32] = 6'h12;
        mem[33] = 6'h17;
        mem[34] = 6'h00;
        mem[35] = 6'h35;
        mem[36] = 6'h1b;
        mem[37] = 6'h06;
        mem[38] = 6'h07;
        mem[39] = 6'h10;
        mem[40] = 6'h3b;
        mem[41] = 6'h3f;
        mem[42] = 6'h0d;
        mem[43] = 6'h3c;
        mem[44] = 6'h08;
        mem[45] = 6'h15;
        mem[46] = 6'h0a;
        mem[47] = 6'h25;
        mem[48] = 6'h03;
        mem[49] = 6'h28;
        mem[50] = 6'h0e;
        mem[51] = 6'h3e;
        mem[52] = 6'h36;
        mem[53] = 6'h3a;
        mem[54] = 6'h2e;
        mem[55] = 6'h21;
        mem[56] = 6'h1d;
        mem[57] = 6'h34;
        mem[58] = 6'h05;
        mem[59] = 6'h0f;
        mem[60] = 6'h01;
        mem[61] = 6'h09;
        mem[62] = 6'h30;
        mem[63] = 6'h0b;
    end
endmodule

module encrypt_4sbox_small8(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h28;
        mem[1] = 6'h3a;
        mem[2] = 6'h30;
        mem[3] = 6'h3f;
        mem[4] = 6'h00;
        mem[5] = 6'h0a;
        mem[6] = 6'h2c;
        mem[7] = 6'h1b;
        mem[8] = 6'h1f;
        mem[9] = 6'h09;
        mem[10] = 6'h38;
        mem[11] = 6'h20;
        mem[12] = 6'h34;
        mem[13] = 6'h2a;
        mem[14] = 6'h2b;
        mem[15] = 6'h15;
        mem[16] = 6'h18;
        mem[17] = 6'h35;
        mem[18] = 6'h21;
        mem[19] = 6'h3d;
        mem[20] = 6'h07;
        mem[21] = 6'h05;
        mem[22] = 6'h10;
        mem[23] = 6'h0f;
        mem[24] = 6'h16;
        mem[25] = 6'h37;
        mem[26] = 6'h2f;
        mem[27] = 6'h0e;
        mem[28] = 6'h23;
        mem[29] = 6'h01;
        mem[30] = 6'h0b;
        mem[31] = 6'h25;
        mem[32] = 6'h31;
        mem[33] = 6'h19;
        mem[34] = 6'h12;
        mem[35] = 6'h2d;
        mem[36] = 6'h1c;
        mem[37] = 6'h3b;
        mem[38] = 6'h03;
        mem[39] = 6'h3e;
        mem[40] = 6'h3c;
        mem[41] = 6'h29;
        mem[42] = 6'h22;
        mem[43] = 6'h13;
        mem[44] = 6'h24;
        mem[45] = 6'h17;
        mem[46] = 6'h1a;
        mem[47] = 6'h02;
        mem[48] = 6'h39;
        mem[49] = 6'h08;
        mem[50] = 6'h26;
        mem[51] = 6'h04;
        mem[52] = 6'h14;
        mem[53] = 6'h32;
        mem[54] = 6'h1e;
        mem[55] = 6'h27;
        mem[56] = 6'h2e;
        mem[57] = 6'h06;
        mem[58] = 6'h33;
        mem[59] = 6'h11;
        mem[60] = 6'h1d;
        mem[61] = 6'h36;
        mem[62] = 6'h0d;
        mem[63] = 6'h0c;
    end
endmodule

module encrypt_4sbox_small9(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h24;
        mem[1] = 6'h1c;
        mem[2] = 6'h0b;
        mem[3] = 6'h2a;
        mem[4] = 6'h0a;
        mem[5] = 6'h36;
        mem[6] = 6'h1a;
        mem[7] = 6'h01;
        mem[8] = 6'h1d;
        mem[9] = 6'h33;
        mem[10] = 6'h3a;
        mem[11] = 6'h37;
        mem[12] = 6'h02;
        mem[13] = 6'h1b;
        mem[14] = 6'h1f;
        mem[15] = 6'h06;
        mem[16] = 6'h07;
        mem[17] = 6'h2d;
        mem[18] = 6'h10;
        mem[19] = 6'h3e;
        mem[20] = 6'h31;
        mem[21] = 6'h39;
        mem[22] = 6'h3b;
        mem[23] = 6'h28;
        mem[24] = 6'h16;
        mem[25] = 6'h23;
        mem[26] = 6'h03;
        mem[27] = 6'h00;
        mem[28] = 6'h0e;
        mem[29] = 6'h2b;
        mem[30] = 6'h0f;
        mem[31] = 6'h29;
        mem[32] = 6'h38;
        mem[33] = 6'h32;
        mem[34] = 6'h19;
        mem[35] = 6'h14;
        mem[36] = 6'h08;
        mem[37] = 6'h09;
        mem[38] = 6'h13;
        mem[39] = 6'h25;
        mem[40] = 6'h3f;
        mem[41] = 6'h35;
        mem[42] = 6'h27;
        mem[43] = 6'h17;
        mem[44] = 6'h30;
        mem[45] = 6'h21;
        mem[46] = 6'h22;
        mem[47] = 6'h3c;
        mem[48] = 6'h1e;
        mem[49] = 6'h0d;
        mem[50] = 6'h18;
        mem[51] = 6'h34;
        mem[52] = 6'h15;
        mem[53] = 6'h3d;
        mem[54] = 6'h11;
        mem[55] = 6'h2f;
        mem[56] = 6'h2e;
        mem[57] = 6'h26;
        mem[58] = 6'h0c;
        mem[59] = 6'h20;
        mem[60] = 6'h05;
        mem[61] = 6'h04;
        mem[62] = 6'h2c;
        mem[63] = 6'h12;
    end
endmodule

module encrypt_4sbox_small10(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h3a;
        mem[1] = 6'h36;
        mem[2] = 6'h2b;
        mem[3] = 6'h1d;
        mem[4] = 6'h03;
        mem[5] = 6'h23;
        mem[6] = 6'h10;
        mem[7] = 6'h3f;
        mem[8] = 6'h2f;
        mem[9] = 6'h22;
        mem[10] = 6'h1f;
        mem[11] = 6'h39;
        mem[12] = 6'h08;
        mem[13] = 6'h32;
        mem[14] = 6'h02;
        mem[15] = 6'h29;
        mem[16] = 6'h14;
        mem[17] = 6'h17;
        mem[18] = 6'h21;
        mem[19] = 6'h20;
        mem[20] = 6'h0c;
        mem[21] = 6'h2c;
        mem[22] = 6'h06;
        mem[23] = 6'h19;
        mem[24] = 6'h3d;
        mem[25] = 6'h11;
        mem[26] = 6'h30;
        mem[27] = 6'h33;
        mem[28] = 6'h16;
        mem[29] = 6'h0e;
        mem[30] = 6'h27;
        mem[31] = 6'h24;
        mem[32] = 6'h26;
        mem[33] = 6'h01;
        mem[34] = 6'h09;
        mem[35] = 6'h25;
        mem[36] = 6'h1a;
        mem[37] = 6'h3b;
        mem[38] = 6'h2e;
        mem[39] = 6'h3e;
        mem[40] = 6'h0f;
        mem[41] = 6'h28;
        mem[42] = 6'h37;
        mem[43] = 6'h2a;
        mem[44] = 6'h35;
        mem[45] = 6'h12;
        mem[46] = 6'h0d;
        mem[47] = 6'h1e;
        mem[48] = 6'h18;
        mem[49] = 6'h04;
        mem[50] = 6'h07;
        mem[51] = 6'h0a;
        mem[52] = 6'h0b;
        mem[53] = 6'h00;
        mem[54] = 6'h3c;
        mem[55] = 6'h31;
        mem[56] = 6'h1b;
        mem[57] = 6'h38;
        mem[58] = 6'h13;
        mem[59] = 6'h2d;
        mem[60] = 6'h15;
        mem[61] = 6'h1c;
        mem[62] = 6'h05;
        mem[63] = 6'h34;
    end
endmodule

module encrypt_4sbox_small11(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h0a;
        mem[1] = 6'h08;
        mem[2] = 6'h1d;
        mem[3] = 6'h2f;
        mem[4] = 6'h06;
        mem[5] = 6'h32;
        mem[6] = 6'h2a;
        mem[7] = 6'h38;
        mem[8] = 6'h37;
        mem[9] = 6'h1f;
        mem[10] = 6'h13;
        mem[11] = 6'h20;
        mem[12] = 6'h11;
        mem[13] = 6'h24;
        mem[14] = 6'h2c;
        mem[15] = 6'h03;
        mem[16] = 6'h36;
        mem[17] = 6'h21;
        mem[18] = 6'h0f;
        mem[19] = 6'h33;
        mem[20] = 6'h1e;
        mem[21] = 6'h1c;
        mem[22] = 6'h0b;
        mem[23] = 6'h28;
        mem[24] = 6'h22;
        mem[25] = 6'h3b;
        mem[26] = 6'h0d;
        mem[27] = 6'h3a;
        mem[28] = 6'h35;
        mem[29] = 6'h2d;
        mem[30] = 6'h07;
        mem[31] = 6'h18;
        mem[32] = 6'h3f;
        mem[33] = 6'h15;
        mem[34] = 6'h25;
        mem[35] = 6'h05;
        mem[36] = 6'h3d;
        mem[37] = 6'h29;
        mem[38] = 6'h02;
        mem[39] = 6'h2b;
        mem[40] = 6'h30;
        mem[41] = 6'h34;
        mem[42] = 6'h10;
        mem[43] = 6'h23;
        mem[44] = 6'h3c;
        mem[45] = 6'h00;
        mem[46] = 6'h16;
        mem[47] = 6'h2e;
        mem[48] = 6'h39;
        mem[49] = 6'h19;
        mem[50] = 6'h1a;
        mem[51] = 6'h1b;
        mem[52] = 6'h27;
        mem[53] = 6'h0e;
        mem[54] = 6'h01;
        mem[55] = 6'h17;
        mem[56] = 6'h26;
        mem[57] = 6'h09;
        mem[58] = 6'h12;
        mem[59] = 6'h0c;
        mem[60] = 6'h3e;
        mem[61] = 6'h14;
        mem[62] = 6'h04;
        mem[63] = 6'h31;
    end
endmodule

module encrypt_4sbox_small12(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h10;
        mem[1] = 6'h3f;
        mem[2] = 6'h15;
        mem[3] = 6'h01;
        mem[4] = 6'h08;
        mem[5] = 6'h1f;
        mem[6] = 6'h23;
        mem[7] = 6'h17;
        mem[8] = 6'h18;
        mem[9] = 6'h02;
        mem[10] = 6'h22;
        mem[11] = 6'h04;
        mem[12] = 6'h33;
        mem[13] = 6'h05;
        mem[14] = 6'h13;
        mem[15] = 6'h3e;
        mem[16] = 6'h2c;
        mem[17] = 6'h0e;
        mem[18] = 6'h27;
        mem[19] = 6'h35;
        mem[20] = 6'h00;
        mem[21] = 6'h39;
        mem[22] = 6'h14;
        mem[23] = 6'h24;
        mem[24] = 6'h1e;
        mem[25] = 6'h3d;
        mem[26] = 6'h2b;
        mem[27] = 6'h1d;
        mem[28] = 6'h20;
        mem[29] = 6'h0c;
        mem[30] = 6'h3a;
        mem[31] = 6'h2d;
        mem[32] = 6'h38;
        mem[33] = 6'h3c;
        mem[34] = 6'h21;
        mem[35] = 6'h29;
        mem[36] = 6'h1c;
        mem[37] = 6'h30;
        mem[38] = 6'h11;
        mem[39] = 6'h0b;
        mem[40] = 6'h36;
        mem[41] = 6'h2f;
        mem[42] = 6'h1b;
        mem[43] = 6'h2a;
        mem[44] = 6'h26;
        mem[45] = 6'h0f;
        mem[46] = 6'h0d;
        mem[47] = 6'h09;
        mem[48] = 6'h34;
        mem[49] = 6'h1a;
        mem[50] = 6'h12;
        mem[51] = 6'h2e;
        mem[52] = 6'h3b;
        mem[53] = 6'h31;
        mem[54] = 6'h03;
        mem[55] = 6'h0a;
        mem[56] = 6'h16;
        mem[57] = 6'h28;
        mem[58] = 6'h19;
        mem[59] = 6'h06;
        mem[60] = 6'h25;
        mem[61] = 6'h07;
        mem[62] = 6'h37;
        mem[63] = 6'h32;
    end
endmodule

module encrypt_4sbox_small13(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h28;
        mem[1] = 6'h36;
        mem[2] = 6'h3d;
        mem[3] = 6'h2e;
        mem[4] = 6'h30;
        mem[5] = 6'h08;
        mem[6] = 6'h1a;
        mem[7] = 6'h35;
        mem[8] = 6'h0c;
        mem[9] = 6'h2f;
        mem[10] = 6'h39;
        mem[11] = 6'h13;
        mem[12] = 6'h27;
        mem[13] = 6'h10;
        mem[14] = 6'h15;
        mem[15] = 6'h29;
        mem[16] = 6'h12;
        mem[17] = 6'h2a;
        mem[18] = 6'h03;
        mem[19] = 6'h00;
        mem[20] = 6'h18;
        mem[21] = 6'h3f;
        mem[22] = 6'h07;
        mem[23] = 6'h0e;
        mem[24] = 6'h31;
        mem[25] = 6'h22;
        mem[26] = 6'h3c;
        mem[27] = 6'h3e;
        mem[28] = 6'h0d;
        mem[29] = 6'h1f;
        mem[30] = 6'h11;
        mem[31] = 6'h23;
        mem[32] = 6'h06;
        mem[33] = 6'h21;
        mem[34] = 6'h2d;
        mem[35] = 6'h1e;
        mem[36] = 6'h34;
        mem[37] = 6'h3a;
        mem[38] = 6'h17;
        mem[39] = 6'h1d;
        mem[40] = 6'h24;
        mem[41] = 6'h0f;
        mem[42] = 6'h26;
        mem[43] = 6'h0a;
        mem[44] = 6'h16;
        mem[45] = 6'h38;
        mem[46] = 6'h02;
        mem[47] = 6'h01;
        mem[48] = 6'h3b;
        mem[49] = 6'h2b;
        mem[50] = 6'h04;
        mem[51] = 6'h33;
        mem[52] = 6'h25;
        mem[53] = 6'h0b;
        mem[54] = 6'h20;
        mem[55] = 6'h19;
        mem[56] = 6'h32;
        mem[57] = 6'h14;
        mem[58] = 6'h1b;
        mem[59] = 6'h1c;
        mem[60] = 6'h37;
        mem[61] = 6'h09;
        mem[62] = 6'h05;
        mem[63] = 6'h2c;
    end
endmodule

module encrypt_4sbox_small14(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h0f;
        mem[1] = 6'h02;
        mem[2] = 6'h38;
        mem[3] = 6'h39;
        mem[4] = 6'h27;
        mem[5] = 6'h2d;
        mem[6] = 6'h1f;
        mem[7] = 6'h21;
        mem[8] = 6'h34;
        mem[9] = 6'h07;
        mem[10] = 6'h1e;
        mem[11] = 6'h32;
        mem[12] = 6'h23;
        mem[13] = 6'h3c;
        mem[14] = 6'h0c;
        mem[15] = 6'h2b;
        mem[16] = 6'h14;
        mem[17] = 6'h2f;
        mem[18] = 6'h16;
        mem[19] = 6'h1c;
        mem[20] = 6'h06;
        mem[21] = 6'h09;
        mem[22] = 6'h20;
        mem[23] = 6'h0e;
        mem[24] = 6'h3f;
        mem[25] = 6'h3d;
        mem[26] = 6'h31;
        mem[27] = 6'h12;
        mem[28] = 6'h1d;
        mem[29] = 6'h25;
        mem[30] = 6'h18;
        mem[31] = 6'h26;
        mem[32] = 6'h2a;
        mem[33] = 6'h0b;
        mem[34] = 6'h35;
        mem[35] = 6'h08;
        mem[36] = 6'h24;
        mem[37] = 6'h05;
        mem[38] = 6'h37;
        mem[39] = 6'h0d;
        mem[40] = 6'h1a;
        mem[41] = 6'h2c;
        mem[42] = 6'h33;
        mem[43] = 6'h3e;
        mem[44] = 6'h29;
        mem[45] = 6'h13;
        mem[46] = 6'h2e;
        mem[47] = 6'h11;
        mem[48] = 6'h15;
        mem[49] = 6'h19;
        mem[50] = 6'h0a;
        mem[51] = 6'h17;
        mem[52] = 6'h03;
        mem[53] = 6'h3b;
        mem[54] = 6'h1b;
        mem[55] = 6'h22;
        mem[56] = 6'h01;
        mem[57] = 6'h00;
        mem[58] = 6'h30;
        mem[59] = 6'h3a;
        mem[60] = 6'h28;
        mem[61] = 6'h10;
        mem[62] = 6'h36;
        mem[63] = 6'h04;
    end
endmodule

module encrypt_4sbox_small15(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h2e;
        mem[1] = 6'h18;
        mem[2] = 6'h11;
        mem[3] = 6'h14;
        mem[4] = 6'h30;
        mem[5] = 6'h23;
        mem[6] = 6'h01;
        mem[7] = 6'h20;
        mem[8] = 6'h2a;
        mem[9] = 6'h1c;
        mem[10] = 6'h27;
        mem[11] = 6'h08;
        mem[12] = 6'h3d;
        mem[13] = 6'h39;
        mem[14] = 6'h04;
        mem[15] = 6'h36;
        mem[16] = 6'h29;
        mem[17] = 6'h3c;
        mem[18] = 6'h32;
        mem[19] = 6'h19;
        mem[20] = 6'h2d;
        mem[21] = 6'h21;
        mem[22] = 6'h3a;
        mem[23] = 6'h35;
        mem[24] = 6'h37;
        mem[25] = 6'h34;
        mem[26] = 6'h0b;
        mem[27] = 6'h03;
        mem[28] = 6'h2f;
        mem[29] = 6'h1a;
        mem[30] = 6'h24;
        mem[31] = 6'h3b;
        mem[32] = 6'h02;
        mem[33] = 6'h2b;
        mem[34] = 6'h0c;
        mem[35] = 6'h06;
        mem[36] = 6'h3e;
        mem[37] = 6'h25;
        mem[38] = 6'h0d;
        mem[39] = 6'h26;
        mem[40] = 6'h09;
        mem[41] = 6'h38;
        mem[42] = 6'h3f;
        mem[43] = 6'h33;
        mem[44] = 6'h31;
        mem[45] = 6'h13;
        mem[46] = 6'h16;
        mem[47] = 6'h1b;
        mem[48] = 6'h1d;
        mem[49] = 6'h17;
        mem[50] = 6'h12;
        mem[51] = 6'h0e;
        mem[52] = 6'h07;
        mem[53] = 6'h0f;
        mem[54] = 6'h10;
        mem[55] = 6'h1f;
        mem[56] = 6'h2c;
        mem[57] = 6'h1e;
        mem[58] = 6'h28;
        mem[59] = 6'h15;
        mem[60] = 6'h0a;
        mem[61] = 6'h05;
        mem[62] = 6'h00;
        mem[63] = 6'h22;
    end
endmodule

module encrypt_4sbox_small16(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h26;
        mem[1] = 6'h2c;
        mem[2] = 6'h0c;
        mem[3] = 6'h2f;
        mem[4] = 6'h0b;
        mem[5] = 6'h0d;
        mem[6] = 6'h18;
        mem[7] = 6'h34;
        mem[8] = 6'h17;
        mem[9] = 6'h30;
        mem[10] = 6'h3d;
        mem[11] = 6'h1c;
        mem[12] = 6'h2b;
        mem[13] = 6'h25;
        mem[14] = 6'h3c;
        mem[15] = 6'h2e;
        mem[16] = 6'h29;
        mem[17] = 6'h36;
        mem[18] = 6'h23;
        mem[19] = 6'h07;
        mem[20] = 6'h14;
        mem[21] = 6'h27;
        mem[22] = 6'h11;
        mem[23] = 6'h08;
        mem[24] = 6'h15;
        mem[25] = 6'h20;
        mem[26] = 6'h3f;
        mem[27] = 6'h22;
        mem[28] = 6'h0e;
        mem[29] = 6'h35;
        mem[30] = 6'h0f;
        mem[31] = 6'h2d;
        mem[32] = 6'h00;
        mem[33] = 6'h19;
        mem[34] = 6'h13;
        mem[35] = 6'h16;
        mem[36] = 6'h12;
        mem[37] = 6'h1d;
        mem[38] = 6'h06;
        mem[39] = 6'h05;
        mem[40] = 6'h1e;
        mem[41] = 6'h09;
        mem[42] = 6'h38;
        mem[43] = 6'h32;
        mem[44] = 6'h28;
        mem[45] = 6'h04;
        mem[46] = 6'h21;
        mem[47] = 6'h1a;
        mem[48] = 6'h3b;
        mem[49] = 6'h37;
        mem[50] = 6'h31;
        mem[51] = 6'h33;
        mem[52] = 6'h02;
        mem[53] = 6'h39;
        mem[54] = 6'h2a;
        mem[55] = 6'h1b;
        mem[56] = 6'h1f;
        mem[57] = 6'h0a;
        mem[58] = 6'h3a;
        mem[59] = 6'h01;
        mem[60] = 6'h3e;
        mem[61] = 6'h24;
        mem[62] = 6'h10;
        mem[63] = 6'h03;
    end
endmodule

module encrypt_4sbox_small17(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h05;
        mem[1] = 6'h34;
        mem[2] = 6'h1a;
        mem[3] = 6'h0d;
        mem[4] = 6'h00;
        mem[5] = 6'h36;
        mem[6] = 6'h02;
        mem[7] = 6'h1f;
        mem[8] = 6'h12;
        mem[9] = 6'h32;
        mem[10] = 6'h2e;
        mem[11] = 6'h3d;
        mem[12] = 6'h3b;
        mem[13] = 6'h33;
        mem[14] = 6'h09;
        mem[15] = 6'h08;
        mem[16] = 6'h06;
        mem[17] = 6'h18;
        mem[18] = 6'h23;
        mem[19] = 6'h1c;
        mem[20] = 6'h16;
        mem[21] = 6'h1b;
        mem[22] = 6'h38;
        mem[23] = 6'h2a;
        mem[24] = 6'h3c;
        mem[25] = 6'h13;
        mem[26] = 6'h3e;
        mem[27] = 6'h22;
        mem[28] = 6'h0b;
        mem[29] = 6'h14;
        mem[30] = 6'h0c;
        mem[31] = 6'h24;
        mem[32] = 6'h25;
        mem[33] = 6'h30;
        mem[34] = 6'h3a;
        mem[35] = 6'h04;
        mem[36] = 6'h10;
        mem[37] = 6'h03;
        mem[38] = 6'h2b;
        mem[39] = 6'h26;
        mem[40] = 6'h31;
        mem[41] = 6'h21;
        mem[42] = 6'h2d;
        mem[43] = 6'h17;
        mem[44] = 6'h3f;
        mem[45] = 6'h35;
        mem[46] = 6'h07;
        mem[47] = 6'h29;
        mem[48] = 6'h37;
        mem[49] = 6'h15;
        mem[50] = 6'h39;
        mem[51] = 6'h2c;
        mem[52] = 6'h0a;
        mem[53] = 6'h28;
        mem[54] = 6'h0f;
        mem[55] = 6'h20;
        mem[56] = 6'h2f;
        mem[57] = 6'h01;
        mem[58] = 6'h11;
        mem[59] = 6'h1d;
        mem[60] = 6'h27;
        mem[61] = 6'h19;
        mem[62] = 6'h1e;
        mem[63] = 6'h0e;
    end
endmodule

module encrypt_4sbox_small18(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h0f;
        mem[1] = 6'h3f;
        mem[2] = 6'h05;
        mem[3] = 6'h17;
        mem[4] = 6'h11;
        mem[5] = 6'h38;
        mem[6] = 6'h1f;
        mem[7] = 6'h14;
        mem[8] = 6'h03;
        mem[9] = 6'h22;
        mem[10] = 6'h37;
        mem[11] = 6'h09;
        mem[12] = 6'h2c;
        mem[13] = 6'h27;
        mem[14] = 6'h1a;
        mem[15] = 6'h19;
        mem[16] = 6'h0d;
        mem[17] = 6'h23;
        mem[18] = 6'h06;
        mem[19] = 6'h25;
        mem[20] = 6'h31;
        mem[21] = 6'h1d;
        mem[22] = 6'h04;
        mem[23] = 6'h29;
        mem[24] = 6'h20;
        mem[25] = 6'h2a;
        mem[26] = 6'h32;
        mem[27] = 6'h0c;
        mem[28] = 6'h3b;
        mem[29] = 6'h39;
        mem[30] = 6'h1c;
        mem[31] = 6'h2b;
        mem[32] = 6'h28;
        mem[33] = 6'h2e;
        mem[34] = 6'h35;
        mem[35] = 6'h3e;
        mem[36] = 6'h10;
        mem[37] = 6'h30;
        mem[38] = 6'h00;
        mem[39] = 6'h1e;
        mem[40] = 6'h34;
        mem[41] = 6'h1b;
        mem[42] = 6'h33;
        mem[43] = 6'h24;
        mem[44] = 6'h2d;
        mem[45] = 6'h12;
        mem[46] = 6'h36;
        mem[47] = 6'h0e;
        mem[48] = 6'h13;
        mem[49] = 6'h0b;
        mem[50] = 6'h3c;
        mem[51] = 6'h2f;
        mem[52] = 6'h15;
        mem[53] = 6'h26;
        mem[54] = 6'h16;
        mem[55] = 6'h3d;
        mem[56] = 6'h21;
        mem[57] = 6'h08;
        mem[58] = 6'h3a;
        mem[59] = 6'h02;
        mem[60] = 6'h0a;
        mem[61] = 6'h18;
        mem[62] = 6'h01;
        mem[63] = 6'h07;
    end
endmodule

module encrypt_4sbox_small19(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h02;
        mem[1] = 6'h11;
        mem[2] = 6'h32;
        mem[3] = 6'h24;
        mem[4] = 6'h0c;
        mem[5] = 6'h33;
        mem[6] = 6'h2f;
        mem[7] = 6'h03;
        mem[8] = 6'h14;
        mem[9] = 6'h3b;
        mem[10] = 6'h1d;
        mem[11] = 6'h0b;
        mem[12] = 6'h35;
        mem[13] = 6'h08;
        mem[14] = 6'h05;
        mem[15] = 6'h06;
        mem[16] = 6'h21;
        mem[17] = 6'h39;
        mem[18] = 6'h36;
        mem[19] = 6'h17;
        mem[20] = 6'h12;
        mem[21] = 6'h38;
        mem[22] = 6'h30;
        mem[23] = 6'h23;
        mem[24] = 6'h19;
        mem[25] = 6'h25;
        mem[26] = 6'h0d;
        mem[27] = 6'h0a;
        mem[28] = 6'h1e;
        mem[29] = 6'h2e;
        mem[30] = 6'h1a;
        mem[31] = 6'h28;
        mem[32] = 6'h1b;
        mem[33] = 6'h2d;
        mem[34] = 6'h20;
        mem[35] = 6'h26;
        mem[36] = 6'h07;
        mem[37] = 6'h2b;
        mem[38] = 6'h34;
        mem[39] = 6'h18;
        mem[40] = 6'h22;
        mem[41] = 6'h1f;
        mem[42] = 6'h2c;
        mem[43] = 6'h01;
        mem[44] = 6'h29;
        mem[45] = 6'h10;
        mem[46] = 6'h3f;
        mem[47] = 6'h0f;
        mem[48] = 6'h3d;
        mem[49] = 6'h16;
        mem[50] = 6'h15;
        mem[51] = 6'h3e;
        mem[52] = 6'h13;
        mem[53] = 6'h37;
        mem[54] = 6'h31;
        mem[55] = 6'h3a;
        mem[56] = 6'h00;
        mem[57] = 6'h3c;
        mem[58] = 6'h1c;
        mem[59] = 6'h27;
        mem[60] = 6'h2a;
        mem[61] = 6'h0e;
        mem[62] = 6'h09;
        mem[63] = 6'h04;
    end
endmodule

module encrypt_4sbox_small20(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h2a;
        mem[1] = 6'h0d;
        mem[2] = 6'h01;
        mem[3] = 6'h13;
        mem[4] = 6'h1a;
        mem[5] = 6'h34;
        mem[6] = 6'h2d;
        mem[7] = 6'h12;
        mem[8] = 6'h23;
        mem[9] = 6'h1b;
        mem[10] = 6'h19;
        mem[11] = 6'h0f;
        mem[12] = 6'h21;
        mem[13] = 6'h09;
        mem[14] = 6'h3b;
        mem[15] = 6'h20;
        mem[16] = 6'h03;
        mem[17] = 6'h1c;
        mem[18] = 6'h24;
        mem[19] = 6'h30;
        mem[20] = 6'h38;
        mem[21] = 6'h32;
        mem[22] = 6'h10;
        mem[23] = 6'h06;
        mem[24] = 6'h35;
        mem[25] = 6'h18;
        mem[26] = 6'h0e;
        mem[27] = 6'h26;
        mem[28] = 6'h1f;
        mem[29] = 6'h27;
        mem[30] = 6'h08;
        mem[31] = 6'h04;
        mem[32] = 6'h3e;
        mem[33] = 6'h15;
        mem[34] = 6'h3d;
        mem[35] = 6'h22;
        mem[36] = 6'h1d;
        mem[37] = 6'h39;
        mem[38] = 6'h2e;
        mem[39] = 6'h1e;
        mem[40] = 6'h37;
        mem[41] = 6'h0b;
        mem[42] = 6'h0c;
        mem[43] = 6'h14;
        mem[44] = 6'h07;
        mem[45] = 6'h3a;
        mem[46] = 6'h33;
        mem[47] = 6'h2c;
        mem[48] = 6'h28;
        mem[49] = 6'h00;
        mem[50] = 6'h2f;
        mem[51] = 6'h11;
        mem[52] = 6'h17;
        mem[53] = 6'h36;
        mem[54] = 6'h2b;
        mem[55] = 6'h31;
        mem[56] = 6'h05;
        mem[57] = 6'h25;
        mem[58] = 6'h16;
        mem[59] = 6'h0a;
        mem[60] = 6'h29;
        mem[61] = 6'h02;
        mem[62] = 6'h3c;
        mem[63] = 6'h3f;
    end
endmodule

module encrypt_4sbox_small21(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h33;
        mem[1] = 6'h30;
        mem[2] = 6'h3a;
        mem[3] = 6'h19;
        mem[4] = 6'h04;
        mem[5] = 6'h0e;
        mem[6] = 6'h1d;
        mem[7] = 6'h3b;
        mem[8] = 6'h0a;
        mem[9] = 6'h0c;
        mem[10] = 6'h22;
        mem[11] = 6'h1f;
        mem[12] = 6'h23;
        mem[13] = 6'h08;
        mem[14] = 6'h28;
        mem[15] = 6'h3c;
        mem[16] = 6'h1b;
        mem[17] = 6'h2c;
        mem[18] = 6'h13;
        mem[19] = 6'h29;
        mem[20] = 6'h3d;
        mem[21] = 6'h20;
        mem[22] = 6'h3f;
        mem[23] = 6'h34;
        mem[24] = 6'h07;
        mem[25] = 6'h2b;
        mem[26] = 6'h21;
        mem[27] = 6'h26;
        mem[28] = 6'h35;
        mem[29] = 6'h27;
        mem[30] = 6'h32;
        mem[31] = 6'h16;
        mem[32] = 6'h02;
        mem[33] = 6'h0b;
        mem[34] = 6'h1a;
        mem[35] = 6'h2a;
        mem[36] = 6'h05;
        mem[37] = 6'h37;
        mem[38] = 6'h06;
        mem[39] = 6'h39;
        mem[40] = 6'h36;
        mem[41] = 6'h11;
        mem[42] = 6'h1e;
        mem[43] = 6'h14;
        mem[44] = 6'h17;
        mem[45] = 6'h0d;
        mem[46] = 6'h03;
        mem[47] = 6'h1c;
        mem[48] = 6'h12;
        mem[49] = 6'h09;
        mem[50] = 6'h10;
        mem[51] = 6'h01;
        mem[52] = 6'h0f;
        mem[53] = 6'h15;
        mem[54] = 6'h24;
        mem[55] = 6'h38;
        mem[56] = 6'h00;
        mem[57] = 6'h2d;
        mem[58] = 6'h18;
        mem[59] = 6'h2e;
        mem[60] = 6'h25;
        mem[61] = 6'h2f;
        mem[62] = 6'h31;
        mem[63] = 6'h3e;
    end
endmodule

module encrypt_4sbox_small22(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h1a;
        mem[1] = 6'h05;
        mem[2] = 6'h38;
        mem[3] = 6'h04;
        mem[4] = 6'h18;
        mem[5] = 6'h13;
        mem[6] = 6'h32;
        mem[7] = 6'h17;
        mem[8] = 6'h1b;
        mem[9] = 6'h31;
        mem[10] = 6'h2e;
        mem[11] = 6'h03;
        mem[12] = 6'h0b;
        mem[13] = 6'h3e;
        mem[14] = 6'h3f;
        mem[15] = 6'h10;
        mem[16] = 6'h09;
        mem[17] = 6'h22;
        mem[18] = 6'h07;
        mem[19] = 6'h2d;
        mem[20] = 6'h2b;
        mem[21] = 6'h36;
        mem[22] = 6'h21;
        mem[23] = 6'h27;
        mem[24] = 6'h19;
        mem[25] = 6'h08;
        mem[26] = 6'h14;
        mem[27] = 6'h15;
        mem[28] = 6'h28;
        mem[29] = 6'h02;
        mem[30] = 6'h3b;
        mem[31] = 6'h2a;
        mem[32] = 6'h3d;
        mem[33] = 6'h34;
        mem[34] = 6'h0e;
        mem[35] = 6'h0c;
        mem[36] = 6'h1f;
        mem[37] = 6'h24;
        mem[38] = 6'h12;
        mem[39] = 6'h0f;
        mem[40] = 6'h1c;
        mem[41] = 6'h2f;
        mem[42] = 6'h2c;
        mem[43] = 6'h06;
        mem[44] = 6'h20;
        mem[45] = 6'h25;
        mem[46] = 6'h35;
        mem[47] = 6'h29;
        mem[48] = 6'h0d;
        mem[49] = 6'h1e;
        mem[50] = 6'h0a;
        mem[51] = 6'h26;
        mem[52] = 6'h30;
        mem[53] = 6'h37;
        mem[54] = 6'h01;
        mem[55] = 6'h11;
        mem[56] = 6'h3c;
        mem[57] = 6'h00;
        mem[58] = 6'h33;
        mem[59] = 6'h1d;
        mem[60] = 6'h3a;
        mem[61] = 6'h16;
        mem[62] = 6'h23;
        mem[63] = 6'h39;
    end
endmodule

module encrypt_4sbox_small23(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h2e;
        mem[1] = 6'h21;
        mem[2] = 6'h3b;
        mem[3] = 6'h01;
        mem[4] = 6'h24;
        mem[5] = 6'h25;
        mem[6] = 6'h0b;
        mem[7] = 6'h36;
        mem[8] = 6'h04;
        mem[9] = 6'h39;
        mem[10] = 6'h07;
        mem[11] = 6'h19;
        mem[12] = 6'h3c;
        mem[13] = 6'h20;
        mem[14] = 6'h0f;
        mem[15] = 6'h2a;
        mem[16] = 6'h33;
        mem[17] = 6'h28;
        mem[18] = 6'h15;
        mem[19] = 6'h34;
        mem[20] = 6'h1e;
        mem[21] = 6'h09;
        mem[22] = 6'h0c;
        mem[23] = 6'h14;
        mem[24] = 6'h1c;
        mem[25] = 6'h2d;
        mem[26] = 6'h1f;
        mem[27] = 6'h3e;
        mem[28] = 6'h10;
        mem[29] = 6'h27;
        mem[30] = 6'h18;
        mem[31] = 6'h2b;
        mem[32] = 6'h26;
        mem[33] = 6'h38;
        mem[34] = 6'h02;
        mem[35] = 6'h11;
        mem[36] = 6'h3a;
        mem[37] = 6'h03;
        mem[38] = 6'h12;
        mem[39] = 6'h2c;
        mem[40] = 6'h30;
        mem[41] = 6'h17;
        mem[42] = 6'h31;
        mem[43] = 6'h3d;
        mem[44] = 6'h32;
        mem[45] = 6'h37;
        mem[46] = 6'h1b;
        mem[47] = 6'h29;
        mem[48] = 6'h2f;
        mem[49] = 6'h0a;
        mem[50] = 6'h16;
        mem[51] = 6'h0d;
        mem[52] = 6'h1d;
        mem[53] = 6'h35;
        mem[54] = 6'h05;
        mem[55] = 6'h22;
        mem[56] = 6'h23;
        mem[57] = 6'h13;
        mem[58] = 6'h08;
        mem[59] = 6'h0e;
        mem[60] = 6'h3f;
        mem[61] = 6'h1a;
        mem[62] = 6'h06;
        mem[63] = 6'h00;
    end
endmodule

module encrypt_4sbox_small24(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h0f;
        mem[1] = 6'h2a;
        mem[2] = 6'h03;
        mem[3] = 6'h37;
        mem[4] = 6'h0a;
        mem[5] = 6'h26;
        mem[6] = 6'h2f;
        mem[7] = 6'h21;
        mem[8] = 6'h10;
        mem[9] = 6'h1b;
        mem[10] = 6'h19;
        mem[11] = 6'h16;
        mem[12] = 6'h1d;
        mem[13] = 6'h17;
        mem[14] = 6'h22;
        mem[15] = 6'h18;
        mem[16] = 6'h39;
        mem[17] = 6'h34;
        mem[18] = 6'h02;
        mem[19] = 6'h09;
        mem[20] = 6'h3e;
        mem[21] = 6'h15;
        mem[22] = 6'h13;
        mem[23] = 6'h38;
        mem[24] = 6'h0d;
        mem[25] = 6'h0c;
        mem[26] = 6'h3f;
        mem[27] = 6'h0b;
        mem[28] = 6'h2b;
        mem[29] = 6'h11;
        mem[30] = 6'h00;
        mem[31] = 6'h28;
        mem[32] = 6'h24;
        mem[33] = 6'h31;
        mem[34] = 6'h25;
        mem[35] = 6'h14;
        mem[36] = 6'h07;
        mem[37] = 6'h3b;
        mem[38] = 6'h29;
        mem[39] = 6'h1a;
        mem[40] = 6'h33;
        mem[41] = 6'h35;
        mem[42] = 6'h1f;
        mem[43] = 6'h3c;
        mem[44] = 6'h05;
        mem[45] = 6'h27;
        mem[46] = 6'h01;
        mem[47] = 6'h1e;
        mem[48] = 6'h12;
        mem[49] = 6'h06;
        mem[50] = 6'h3d;
        mem[51] = 6'h1c;
        mem[52] = 6'h04;
        mem[53] = 6'h2e;
        mem[54] = 6'h30;
        mem[55] = 6'h3a;
        mem[56] = 6'h08;
        mem[57] = 6'h20;
        mem[58] = 6'h2d;
        mem[59] = 6'h2c;
        mem[60] = 6'h0e;
        mem[61] = 6'h36;
        mem[62] = 6'h32;
        mem[63] = 6'h23;
    end
endmodule

module encrypt_4sbox_small25(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h03;
        mem[1] = 6'h32;
        mem[2] = 6'h07;
        mem[3] = 6'h10;
        mem[4] = 6'h17;
        mem[5] = 6'h20;
        mem[6] = 6'h24;
        mem[7] = 6'h15;
        mem[8] = 6'h36;
        mem[9] = 6'h08;
        mem[10] = 6'h3a;
        mem[11] = 6'h21;
        mem[12] = 6'h00;
        mem[13] = 6'h31;
        mem[14] = 6'h37;
        mem[15] = 6'h13;
        mem[16] = 6'h06;
        mem[17] = 6'h1f;
        mem[18] = 6'h14;
        mem[19] = 6'h2a;
        mem[20] = 6'h2e;
        mem[21] = 6'h11;
        mem[22] = 6'h29;
        mem[23] = 6'h22;
        mem[24] = 6'h01;
        mem[25] = 6'h18;
        mem[26] = 6'h34;
        mem[27] = 6'h30;
        mem[28] = 6'h0a;
        mem[29] = 6'h09;
        mem[30] = 6'h2b;
        mem[31] = 6'h16;
        mem[32] = 6'h1e;
        mem[33] = 6'h3b;
        mem[34] = 6'h2c;
        mem[35] = 6'h25;
        mem[36] = 6'h0c;
        mem[37] = 6'h33;
        mem[38] = 6'h1b;
        mem[39] = 6'h26;
        mem[40] = 6'h38;
        mem[41] = 6'h0b;
        mem[42] = 6'h3d;
        mem[43] = 6'h3f;
        mem[44] = 6'h0e;
        mem[45] = 6'h05;
        mem[46] = 6'h1a;
        mem[47] = 6'h35;
        mem[48] = 6'h39;
        mem[49] = 6'h0f;
        mem[50] = 6'h27;
        mem[51] = 6'h0d;
        mem[52] = 6'h3e;
        mem[53] = 6'h2f;
        mem[54] = 6'h23;
        mem[55] = 6'h1d;
        mem[56] = 6'h12;
        mem[57] = 6'h28;
        mem[58] = 6'h19;
        mem[59] = 6'h02;
        mem[60] = 6'h2d;
        mem[61] = 6'h3c;
        mem[62] = 6'h04;
        mem[63] = 6'h1c;
    end
endmodule

module encrypt_4sbox_small26(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h20;
        mem[1] = 6'h28;
        mem[2] = 6'h1d;
        mem[3] = 6'h3f;
        mem[4] = 6'h11;
        mem[5] = 6'h13;
        mem[6] = 6'h34;
        mem[7] = 6'h2a;
        mem[8] = 6'h02;
        mem[9] = 6'h3b;
        mem[10] = 6'h0e;
        mem[11] = 6'h0c;
        mem[12] = 6'h37;
        mem[13] = 6'h1a;
        mem[14] = 6'h3a;
        mem[15] = 6'h30;
        mem[16] = 6'h05;
        mem[17] = 6'h32;
        mem[18] = 6'h14;
        mem[19] = 6'h10;
        mem[20] = 6'h15;
        mem[21] = 6'h1e;
        mem[22] = 6'h0a;
        mem[23] = 6'h3d;
        mem[24] = 6'h25;
        mem[25] = 6'h01;
        mem[26] = 6'h1b;
        mem[27] = 6'h24;
        mem[28] = 6'h31;
        mem[29] = 6'h12;
        mem[30] = 6'h07;
        mem[31] = 6'h2d;
        mem[32] = 6'h35;
        mem[33] = 6'h29;
        mem[34] = 6'h03;
        mem[35] = 6'h26;
        mem[36] = 6'h38;
        mem[37] = 6'h18;
        mem[38] = 6'h39;
        mem[39] = 6'h36;
        mem[40] = 6'h00;
        mem[41] = 6'h27;
        mem[42] = 6'h3c;
        mem[43] = 6'h1f;
        mem[44] = 6'h2f;
        mem[45] = 6'h2e;
        mem[46] = 6'h33;
        mem[47] = 6'h0f;
        mem[48] = 6'h2c;
        mem[49] = 6'h06;
        mem[50] = 6'h0d;
        mem[51] = 6'h1c;
        mem[52] = 6'h3e;
        mem[53] = 6'h16;
        mem[54] = 6'h0b;
        mem[55] = 6'h09;
        mem[56] = 6'h23;
        mem[57] = 6'h2b;
        mem[58] = 6'h04;
        mem[59] = 6'h19;
        mem[60] = 6'h21;
        mem[61] = 6'h17;
        mem[62] = 6'h22;
        mem[63] = 6'h08;
    end
endmodule

module encrypt_4sbox_small27(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h25;
        mem[1] = 6'h12;
        mem[2] = 6'h1a;
        mem[3] = 6'h0b;
        mem[4] = 6'h21;
        mem[5] = 6'h1b;
        mem[6] = 6'h36;
        mem[7] = 6'h03;
        mem[8] = 6'h35;
        mem[9] = 6'h14;
        mem[10] = 6'h08;
        mem[11] = 6'h0e;
        mem[12] = 6'h28;
        mem[13] = 6'h39;
        mem[14] = 6'h27;
        mem[15] = 6'h11;
        mem[16] = 6'h0a;
        mem[17] = 6'h16;
        mem[18] = 6'h04;
        mem[19] = 6'h0c;
        mem[20] = 6'h06;
        mem[21] = 6'h2d;
        mem[22] = 6'h22;
        mem[23] = 6'h37;
        mem[24] = 6'h2e;
        mem[25] = 6'h3b;
        mem[26] = 6'h2f;
        mem[27] = 6'h01;
        mem[28] = 6'h1d;
        mem[29] = 6'h1e;
        mem[30] = 6'h17;
        mem[31] = 6'h3c;
        mem[32] = 6'h29;
        mem[33] = 6'h38;
        mem[34] = 6'h24;
        mem[35] = 6'h18;
        mem[36] = 6'h26;
        mem[37] = 6'h3f;
        mem[38] = 6'h07;
        mem[39] = 6'h23;
        mem[40] = 6'h13;
        mem[41] = 6'h2c;
        mem[42] = 6'h3d;
        mem[43] = 6'h32;
        mem[44] = 6'h2a;
        mem[45] = 6'h00;
        mem[46] = 6'h15;
        mem[47] = 6'h05;
        mem[48] = 6'h20;
        mem[49] = 6'h3a;
        mem[50] = 6'h0f;
        mem[51] = 6'h1c;
        mem[52] = 6'h2b;
        mem[53] = 6'h10;
        mem[54] = 6'h31;
        mem[55] = 6'h0d;
        mem[56] = 6'h30;
        mem[57] = 6'h1f;
        mem[58] = 6'h09;
        mem[59] = 6'h02;
        mem[60] = 6'h19;
        mem[61] = 6'h33;
        mem[62] = 6'h34;
        mem[63] = 6'h3e;
    end
endmodule

module encrypt_4sbox_small28(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h08;
        mem[1] = 6'h31;
        mem[2] = 6'h37;
        mem[3] = 6'h1c;
        mem[4] = 6'h25;
        mem[5] = 6'h26;
        mem[6] = 6'h13;
        mem[7] = 6'h0f;
        mem[8] = 6'h10;
        mem[9] = 6'h03;
        mem[10] = 6'h2a;
        mem[11] = 6'h15;
        mem[12] = 6'h30;
        mem[13] = 6'h29;
        mem[14] = 6'h09;
        mem[15] = 6'h28;
        mem[16] = 6'h18;
        mem[17] = 6'h3f;
        mem[18] = 6'h01;
        mem[19] = 6'h23;
        mem[20] = 6'h02;
        mem[21] = 6'h0c;
        mem[22] = 6'h32;
        mem[23] = 6'h36;
        mem[24] = 6'h1e;
        mem[25] = 6'h3d;
        mem[26] = 6'h2d;
        mem[27] = 6'h17;
        mem[28] = 6'h3e;
        mem[29] = 6'h0a;
        mem[30] = 6'h20;
        mem[31] = 6'h12;
        mem[32] = 6'h27;
        mem[33] = 6'h2e;
        mem[34] = 6'h14;
        mem[35] = 6'h35;
        mem[36] = 6'h0d;
        mem[37] = 6'h2f;
        mem[38] = 6'h06;
        mem[39] = 6'h16;
        mem[40] = 6'h3a;
        mem[41] = 6'h3b;
        mem[42] = 6'h33;
        mem[43] = 6'h11;
        mem[44] = 6'h00;
        mem[45] = 6'h04;
        mem[46] = 6'h2b;
        mem[47] = 6'h22;
        mem[48] = 6'h1b;
        mem[49] = 6'h1d;
        mem[50] = 6'h0e;
        mem[51] = 6'h0b;
        mem[52] = 6'h38;
        mem[53] = 6'h19;
        mem[54] = 6'h24;
        mem[55] = 6'h39;
        mem[56] = 6'h21;
        mem[57] = 6'h05;
        mem[58] = 6'h34;
        mem[59] = 6'h1a;
        mem[60] = 6'h2c;
        mem[61] = 6'h3c;
        mem[62] = 6'h1f;
        mem[63] = 6'h07;
    end
endmodule

module encrypt_4sbox_small29(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h2b;
        mem[1] = 6'h3c;
        mem[2] = 6'h29;
        mem[3] = 6'h20;
        mem[4] = 6'h17;
        mem[5] = 6'h14;
        mem[6] = 6'h28;
        mem[7] = 6'h04;
        mem[8] = 6'h21;
        mem[9] = 6'h30;
        mem[10] = 6'h3b;
        mem[11] = 6'h2e;
        mem[12] = 6'h25;
        mem[13] = 6'h37;
        mem[14] = 6'h02;
        mem[15] = 6'h16;
        mem[16] = 6'h12;
        mem[17] = 6'h11;
        mem[18] = 6'h0b;
        mem[19] = 6'h2f;
        mem[20] = 6'h34;
        mem[21] = 6'h3d;
        mem[22] = 6'h0c;
        mem[23] = 6'h2c;
        mem[24] = 6'h1b;
        mem[25] = 6'h3f;
        mem[26] = 6'h31;
        mem[27] = 6'h27;
        mem[28] = 6'h23;
        mem[29] = 6'h01;
        mem[30] = 6'h13;
        mem[31] = 6'h0f;
        mem[32] = 6'h33;
        mem[33] = 6'h1f;
        mem[34] = 6'h3e;
        mem[35] = 6'h2a;
        mem[36] = 6'h24;
        mem[37] = 6'h0a;
        mem[38] = 6'h3a;
        mem[39] = 6'h32;
        mem[40] = 6'h2d;
        mem[41] = 6'h09;
        mem[42] = 6'h19;
        mem[43] = 6'h1e;
        mem[44] = 6'h39;
        mem[45] = 6'h0e;
        mem[46] = 6'h35;
        mem[47] = 6'h26;
        mem[48] = 6'h18;
        mem[49] = 6'h06;
        mem[50] = 6'h05;
        mem[51] = 6'h03;
        mem[52] = 6'h15;
        mem[53] = 6'h38;
        mem[54] = 6'h36;
        mem[55] = 6'h1c;
        mem[56] = 6'h00;
        mem[57] = 6'h08;
        mem[58] = 6'h07;
        mem[59] = 6'h1a;
        mem[60] = 6'h22;
        mem[61] = 6'h1d;
        mem[62] = 6'h10;
        mem[63] = 6'h0d;
    end
endmodule

module encrypt_4sbox_small30(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h12;
        mem[1] = 6'h0a;
        mem[2] = 6'h38;
        mem[3] = 6'h25;
        mem[4] = 6'h02;
        mem[5] = 6'h2e;
        mem[6] = 6'h1e;
        mem[7] = 6'h21;
        mem[8] = 6'h32;
        mem[9] = 6'h1c;
        mem[10] = 6'h1d;
        mem[11] = 6'h3b;
        mem[12] = 6'h04;
        mem[13] = 6'h09;
        mem[14] = 6'h18;
        mem[15] = 6'h3e;
        mem[16] = 6'h31;
        mem[17] = 6'h3d;
        mem[18] = 6'h3c;
        mem[19] = 6'h2c;
        mem[20] = 6'h34;
        mem[21] = 6'h35;
        mem[22] = 6'h14;
        mem[23] = 6'h13;
        mem[24] = 6'h11;
        mem[25] = 6'h22;
        mem[26] = 6'h26;
        mem[27] = 6'h33;
        mem[28] = 6'h24;
        mem[29] = 6'h16;
        mem[30] = 6'h30;
        mem[31] = 6'h3f;
        mem[32] = 6'h2b;
        mem[33] = 6'h2a;
        mem[34] = 6'h23;
        mem[35] = 6'h03;
        mem[36] = 6'h0f;
        mem[37] = 6'h00;
        mem[38] = 6'h2f;
        mem[39] = 6'h27;
        mem[40] = 6'h36;
        mem[41] = 6'h06;
        mem[42] = 6'h15;
        mem[43] = 6'h1b;
        mem[44] = 6'h28;
        mem[45] = 6'h20;
        mem[46] = 6'h05;
        mem[47] = 6'h1f;
        mem[48] = 6'h01;
        mem[49] = 6'h19;
        mem[50] = 6'h39;
        mem[51] = 6'h0d;
        mem[52] = 6'h29;
        mem[53] = 6'h0c;
        mem[54] = 6'h07;
        mem[55] = 6'h17;
        mem[56] = 6'h2d;
        mem[57] = 6'h0e;
        mem[58] = 6'h08;
        mem[59] = 6'h10;
        mem[60] = 6'h3a;
        mem[61] = 6'h0b;
        mem[62] = 6'h1a;
        mem[63] = 6'h37;
    end
endmodule

module encrypt_4sbox_small31(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h3d;
        mem[1] = 6'h0d;
        mem[2] = 6'h34;
        mem[3] = 6'h18;
        mem[4] = 6'h2e;
        mem[5] = 6'h12;
        mem[6] = 6'h14;
        mem[7] = 6'h39;
        mem[8] = 6'h3a;
        mem[9] = 6'h33;
        mem[10] = 6'h10;
        mem[11] = 6'h29;
        mem[12] = 6'h13;
        mem[13] = 6'h30;
        mem[14] = 6'h1c;
        mem[15] = 6'h00;
        mem[16] = 6'h27;
        mem[17] = 6'h28;
        mem[18] = 6'h04;
        mem[19] = 6'h0a;
        mem[20] = 6'h08;
        mem[21] = 6'h0f;
        mem[22] = 6'h3c;
        mem[23] = 6'h24;
        mem[24] = 6'h1a;
        mem[25] = 6'h03;
        mem[26] = 6'h3f;
        mem[27] = 6'h11;
        mem[28] = 6'h25;
        mem[29] = 6'h1d;
        mem[30] = 6'h16;
        mem[31] = 6'h02;
        mem[32] = 6'h38;
        mem[33] = 6'h2f;
        mem[34] = 6'h09;
        mem[35] = 6'h31;
        mem[36] = 6'h2d;
        mem[37] = 6'h15;
        mem[38] = 6'h22;
        mem[39] = 6'h20;
        mem[40] = 6'h32;
        mem[41] = 6'h23;
        mem[42] = 6'h06;
        mem[43] = 6'h2a;
        mem[44] = 6'h01;
        mem[45] = 6'h0c;
        mem[46] = 6'h0e;
        mem[47] = 6'h21;
        mem[48] = 6'h2c;
        mem[49] = 6'h26;
        mem[50] = 6'h3e;
        mem[51] = 6'h0b;
        mem[52] = 6'h1e;
        mem[53] = 6'h35;
        mem[54] = 6'h2b;
        mem[55] = 6'h1f;
        mem[56] = 6'h05;
        mem[57] = 6'h1b;
        mem[58] = 6'h36;
        mem[59] = 6'h07;
        mem[60] = 6'h19;
        mem[61] = 6'h3b;
        mem[62] = 6'h17;
        mem[63] = 6'h37;
    end
endmodule

module encrypt_4sbox_small32(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h0d;
        mem[1] = 6'h00;
        mem[2] = 6'h35;
        mem[3] = 6'h1e;
        mem[4] = 6'h22;
        mem[5] = 6'h20;
        mem[6] = 6'h24;
        mem[7] = 6'h34;
        mem[8] = 6'h18;
        mem[9] = 6'h26;
        mem[10] = 6'h37;
        mem[11] = 6'h1f;
        mem[12] = 6'h1c;
        mem[13] = 6'h10;
        mem[14] = 6'h15;
        mem[15] = 6'h0f;
        mem[16] = 6'h30;
        mem[17] = 6'h31;
        mem[18] = 6'h3a;
        mem[19] = 6'h11;
        mem[20] = 6'h25;
        mem[21] = 6'h36;
        mem[22] = 6'h27;
        mem[23] = 6'h21;
        mem[24] = 6'h1b;
        mem[25] = 6'h3b;
        mem[26] = 6'h1a;
        mem[27] = 6'h28;
        mem[28] = 6'h23;
        mem[29] = 6'h3d;
        mem[30] = 6'h17;
        mem[31] = 6'h29;
        mem[32] = 6'h33;
        mem[33] = 6'h05;
        mem[34] = 6'h0a;
        mem[35] = 6'h3c;
        mem[36] = 6'h2c;
        mem[37] = 6'h32;
        mem[38] = 6'h02;
        mem[39] = 6'h0c;
        mem[40] = 6'h13;
        mem[41] = 6'h39;
        mem[42] = 6'h2e;
        mem[43] = 6'h12;
        mem[44] = 6'h08;
        mem[45] = 6'h03;
        mem[46] = 6'h3f;
        mem[47] = 6'h14;
        mem[48] = 6'h1d;
        mem[49] = 6'h38;
        mem[50] = 6'h04;
        mem[51] = 6'h2b;
        mem[52] = 6'h07;
        mem[53] = 6'h0b;
        mem[54] = 6'h09;
        mem[55] = 6'h3e;
        mem[56] = 6'h19;
        mem[57] = 6'h01;
        mem[58] = 6'h2d;
        mem[59] = 6'h2a;
        mem[60] = 6'h16;
        mem[61] = 6'h0e;
        mem[62] = 6'h2f;
        mem[63] = 6'h06;
    end
endmodule

module encrypt_4sbox_small33(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h35;
        mem[1] = 6'h20;
        mem[2] = 6'h3a;
        mem[3] = 6'h2c;
        mem[4] = 6'h17;
        mem[5] = 6'h27;
        mem[6] = 6'h2f;
        mem[7] = 6'h2b;
        mem[8] = 6'h2e;
        mem[9] = 6'h32;
        mem[10] = 6'h04;
        mem[11] = 6'h22;
        mem[12] = 6'h1c;
        mem[13] = 6'h38;
        mem[14] = 6'h14;
        mem[15] = 6'h0b;
        mem[16] = 6'h26;
        mem[17] = 6'h0e;
        mem[18] = 6'h12;
        mem[19] = 6'h36;
        mem[20] = 6'h05;
        mem[21] = 6'h28;
        mem[22] = 6'h23;
        mem[23] = 6'h39;
        mem[24] = 6'h09;
        mem[25] = 6'h01;
        mem[26] = 6'h0a;
        mem[27] = 6'h1e;
        mem[28] = 6'h13;
        mem[29] = 6'h08;
        mem[30] = 6'h25;
        mem[31] = 6'h34;
        mem[32] = 6'h30;
        mem[33] = 6'h3e;
        mem[34] = 6'h11;
        mem[35] = 6'h21;
        mem[36] = 6'h24;
        mem[37] = 6'h3b;
        mem[38] = 6'h0f;
        mem[39] = 6'h33;
        mem[40] = 6'h31;
        mem[41] = 6'h2d;
        mem[42] = 6'h18;
        mem[43] = 6'h3c;
        mem[44] = 6'h06;
        mem[45] = 6'h29;
        mem[46] = 6'h3f;
        mem[47] = 6'h00;
        mem[48] = 6'h07;
        mem[49] = 6'h02;
        mem[50] = 6'h1d;
        mem[51] = 6'h37;
        mem[52] = 6'h10;
        mem[53] = 6'h15;
        mem[54] = 6'h03;
        mem[55] = 6'h19;
        mem[56] = 6'h16;
        mem[57] = 6'h1f;
        mem[58] = 6'h1b;
        mem[59] = 6'h2a;
        mem[60] = 6'h0d;
        mem[61] = 6'h3d;
        mem[62] = 6'h0c;
        mem[63] = 6'h1a;
    end
endmodule

module encrypt_4sbox_small34(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h2a;
        mem[1] = 6'h37;
        mem[2] = 6'h28;
        mem[3] = 6'h21;
        mem[4] = 6'h2e;
        mem[5] = 6'h22;
        mem[6] = 6'h09;
        mem[7] = 6'h08;
        mem[8] = 6'h39;
        mem[9] = 6'h29;
        mem[10] = 6'h0c;
        mem[11] = 6'h35;
        mem[12] = 6'h3b;
        mem[13] = 6'h14;
        mem[14] = 6'h05;
        mem[15] = 6'h1e;
        mem[16] = 6'h0e;
        mem[17] = 6'h02;
        mem[18] = 6'h27;
        mem[19] = 6'h25;
        mem[20] = 6'h32;
        mem[21] = 6'h20;
        mem[22] = 6'h16;
        mem[23] = 6'h0d;
        mem[24] = 6'h31;
        mem[25] = 6'h07;
        mem[26] = 6'h3f;
        mem[27] = 6'h1a;
        mem[28] = 6'h0f;
        mem[29] = 6'h0a;
        mem[30] = 6'h30;
        mem[31] = 6'h10;
        mem[32] = 6'h23;
        mem[33] = 6'h06;
        mem[34] = 6'h2c;
        mem[35] = 6'h17;
        mem[36] = 6'h11;
        mem[37] = 6'h00;
        mem[38] = 6'h1c;
        mem[39] = 6'h3d;
        mem[40] = 6'h33;
        mem[41] = 6'h15;
        mem[42] = 6'h2d;
        mem[43] = 6'h03;
        mem[44] = 6'h3e;
        mem[45] = 6'h1b;
        mem[46] = 6'h38;
        mem[47] = 6'h26;
        mem[48] = 6'h3a;
        mem[49] = 6'h12;
        mem[50] = 6'h18;
        mem[51] = 6'h19;
        mem[52] = 6'h04;
        mem[53] = 6'h3c;
        mem[54] = 6'h34;
        mem[55] = 6'h1f;
        mem[56] = 6'h13;
        mem[57] = 6'h2f;
        mem[58] = 6'h01;
        mem[59] = 6'h2b;
        mem[60] = 6'h0b;
        mem[61] = 6'h1d;
        mem[62] = 6'h24;
        mem[63] = 6'h36;
    end
endmodule

module encrypt_4sbox_small35(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h3a;
        mem[1] = 6'h1b;
        mem[2] = 6'h02;
        mem[3] = 6'h07;
        mem[4] = 6'h38;
        mem[5] = 6'h37;
        mem[6] = 6'h0a;
        mem[7] = 6'h09;
        mem[8] = 6'h19;
        mem[9] = 6'h20;
        mem[10] = 6'h00;
        mem[11] = 6'h16;
        mem[12] = 6'h1c;
        mem[13] = 6'h1a;
        mem[14] = 6'h23;
        mem[15] = 6'h3c;
        mem[16] = 6'h34;
        mem[17] = 6'h33;
        mem[18] = 6'h2b;
        mem[19] = 6'h35;
        mem[20] = 6'h39;
        mem[21] = 6'h27;
        mem[22] = 6'h28;
        mem[23] = 6'h0b;
        mem[24] = 6'h3e;
        mem[25] = 6'h13;
        mem[26] = 6'h3b;
        mem[27] = 6'h03;
        mem[28] = 6'h2f;
        mem[29] = 6'h05;
        mem[30] = 6'h10;
        mem[31] = 6'h15;
        mem[32] = 6'h1d;
        mem[33] = 6'h14;
        mem[34] = 6'h1f;
        mem[35] = 6'h0d;
        mem[36] = 6'h36;
        mem[37] = 6'h3f;
        mem[38] = 6'h24;
        mem[39] = 6'h01;
        mem[40] = 6'h0e;
        mem[41] = 6'h06;
        mem[42] = 6'h22;
        mem[43] = 6'h26;
        mem[44] = 6'h29;
        mem[45] = 6'h0f;
        mem[46] = 6'h21;
        mem[47] = 6'h31;
        mem[48] = 6'h08;
        mem[49] = 6'h11;
        mem[50] = 6'h1e;
        mem[51] = 6'h3d;
        mem[52] = 6'h17;
        mem[53] = 6'h2d;
        mem[54] = 6'h30;
        mem[55] = 6'h04;
        mem[56] = 6'h25;
        mem[57] = 6'h12;
        mem[58] = 6'h2e;
        mem[59] = 6'h0c;
        mem[60] = 6'h32;
        mem[61] = 6'h18;
        mem[62] = 6'h2c;
        mem[63] = 6'h2a;
    end
endmodule

module encrypt_4sbox_small36(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h11;
        mem[1] = 6'h2f;
        mem[2] = 6'h1f;
        mem[3] = 6'h08;
        mem[4] = 6'h38;
        mem[5] = 6'h16;
        mem[6] = 6'h2e;
        mem[7] = 6'h39;
        mem[8] = 6'h2b;
        mem[9] = 6'h1e;
        mem[10] = 6'h28;
        mem[11] = 6'h00;
        mem[12] = 6'h1d;
        mem[13] = 6'h0a;
        mem[14] = 6'h30;
        mem[15] = 6'h26;
        mem[16] = 6'h32;
        mem[17] = 6'h19;
        mem[18] = 6'h27;
        mem[19] = 6'h3a;
        mem[20] = 6'h35;
        mem[21] = 6'h2d;
        mem[22] = 6'h3c;
        mem[23] = 6'h2a;
        mem[24] = 6'h13;
        mem[25] = 6'h12;
        mem[26] = 6'h01;
        mem[27] = 6'h37;
        mem[28] = 6'h3f;
        mem[29] = 6'h0c;
        mem[30] = 6'h15;
        mem[31] = 6'h34;
        mem[32] = 6'h0f;
        mem[33] = 6'h3e;
        mem[34] = 6'h1c;
        mem[35] = 6'h04;
        mem[36] = 6'h31;
        mem[37] = 6'h29;
        mem[38] = 6'h0e;
        mem[39] = 6'h06;
        mem[40] = 6'h21;
        mem[41] = 6'h17;
        mem[42] = 6'h03;
        mem[43] = 6'h25;
        mem[44] = 6'h36;
        mem[45] = 6'h20;
        mem[46] = 6'h18;
        mem[47] = 6'h14;
        mem[48] = 6'h07;
        mem[49] = 6'h02;
        mem[50] = 6'h22;
        mem[51] = 6'h3d;
        mem[52] = 6'h1b;
        mem[53] = 6'h23;
        mem[54] = 6'h33;
        mem[55] = 6'h0b;
        mem[56] = 6'h3b;
        mem[57] = 6'h0d;
        mem[58] = 6'h05;
        mem[59] = 6'h10;
        mem[60] = 6'h2c;
        mem[61] = 6'h09;
        mem[62] = 6'h24;
        mem[63] = 6'h1a;
    end
endmodule

module encrypt_4sbox_small37(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h00;
        mem[1] = 6'h06;
        mem[2] = 6'h24;
        mem[3] = 6'h02;
        mem[4] = 6'h3d;
        mem[5] = 6'h2d;
        mem[6] = 6'h3c;
        mem[7] = 6'h28;
        mem[8] = 6'h2b;
        mem[9] = 6'h25;
        mem[10] = 6'h16;
        mem[11] = 6'h31;
        mem[12] = 6'h0a;
        mem[13] = 6'h14;
        mem[14] = 6'h17;
        mem[15] = 6'h39;
        mem[16] = 6'h01;
        mem[17] = 6'h20;
        mem[18] = 6'h2a;
        mem[19] = 6'h22;
        mem[20] = 6'h03;
        mem[21] = 6'h2f;
        mem[22] = 6'h30;
        mem[23] = 6'h38;
        mem[24] = 6'h0d;
        mem[25] = 6'h13;
        mem[26] = 6'h04;
        mem[27] = 6'h21;
        mem[28] = 6'h0f;
        mem[29] = 6'h15;
        mem[30] = 6'h33;
        mem[31] = 6'h26;
        mem[32] = 6'h2c;
        mem[33] = 6'h35;
        mem[34] = 6'h12;
        mem[35] = 6'h1f;
        mem[36] = 6'h1e;
        mem[37] = 6'h0b;
        mem[38] = 6'h32;
        mem[39] = 6'h3f;
        mem[40] = 6'h2e;
        mem[41] = 6'h0e;
        mem[42] = 6'h27;
        mem[43] = 6'h1a;
        mem[44] = 6'h37;
        mem[45] = 6'h0c;
        mem[46] = 6'h3e;
        mem[47] = 6'h18;
        mem[48] = 6'h08;
        mem[49] = 6'h10;
        mem[50] = 6'h34;
        mem[51] = 6'h36;
        mem[52] = 6'h29;
        mem[53] = 6'h1b;
        mem[54] = 6'h07;
        mem[55] = 6'h1d;
        mem[56] = 6'h23;
        mem[57] = 6'h09;
        mem[58] = 6'h19;
        mem[59] = 6'h3a;
        mem[60] = 6'h11;
        mem[61] = 6'h05;
        mem[62] = 6'h3b;
        mem[63] = 6'h1c;
    end
endmodule

module encrypt_4sbox_small38(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h07;
        mem[1] = 6'h0d;
        mem[2] = 6'h2f;
        mem[3] = 6'h23;
        mem[4] = 6'h26;
        mem[5] = 6'h09;
        mem[6] = 6'h0e;
        mem[7] = 6'h15;
        mem[8] = 6'h03;
        mem[9] = 6'h20;
        mem[10] = 6'h30;
        mem[11] = 6'h3b;
        mem[12] = 6'h2c;
        mem[13] = 6'h05;
        mem[14] = 6'h16;
        mem[15] = 6'h18;
        mem[16] = 6'h3c;
        mem[17] = 6'h2a;
        mem[18] = 6'h36;
        mem[19] = 6'h3f;
        mem[20] = 6'h38;
        mem[21] = 6'h2d;
        mem[22] = 6'h24;
        mem[23] = 6'h12;
        mem[24] = 6'h1f;
        mem[25] = 6'h3d;
        mem[26] = 6'h1a;
        mem[27] = 6'h39;
        mem[28] = 6'h21;
        mem[29] = 6'h1b;
        mem[30] = 6'h1e;
        mem[31] = 6'h0b;
        mem[32] = 6'h28;
        mem[33] = 6'h10;
        mem[34] = 6'h08;
        mem[35] = 6'h19;
        mem[36] = 6'h33;
        mem[37] = 6'h0f;
        mem[38] = 6'h00;
        mem[39] = 6'h04;
        mem[40] = 6'h27;
        mem[41] = 6'h01;
        mem[42] = 6'h2b;
        mem[43] = 6'h1d;
        mem[44] = 6'h22;
        mem[45] = 6'h29;
        mem[46] = 6'h13;
        mem[47] = 6'h32;
        mem[48] = 6'h25;
        mem[49] = 6'h17;
        mem[50] = 6'h2e;
        mem[51] = 6'h34;
        mem[52] = 6'h3e;
        mem[53] = 6'h1c;
        mem[54] = 6'h02;
        mem[55] = 6'h14;
        mem[56] = 6'h06;
        mem[57] = 6'h37;
        mem[58] = 6'h35;
        mem[59] = 6'h11;
        mem[60] = 6'h3a;
        mem[61] = 6'h0a;
        mem[62] = 6'h0c;
        mem[63] = 6'h31;
    end
endmodule

module encrypt_4sbox_small39(clk, in, out);
    input clk;
    input [5:0] in;
    output reg [5:0] out;
    reg [5:0] mem[0:63];
    always @(posedge clk) begin
        out <= mem[in];
    end
    initial begin
        mem[0] = 6'h17;
        mem[1] = 6'h32;
        mem[2] = 6'h06;
        mem[3] = 6'h2f;
        mem[4] = 6'h28;
        mem[5] = 6'h38;
        mem[6] = 6'h18;
        mem[7] = 6'h26;
        mem[8] = 6'h25;
        mem[9] = 6'h00;
        mem[10] = 6'h27;
        mem[11] = 6'h12;
        mem[12] = 6'h14;
        mem[13] = 6'h29;
        mem[14] = 6'h1d;
        mem[15] = 6'h35;
        mem[16] = 6'h08;
        mem[17] = 6'h3e;
        mem[18] = 6'h0d;
        mem[19] = 6'h34;
        mem[20] = 6'h37;
        mem[21] = 6'h07;
        mem[22] = 6'h1e;
        mem[23] = 6'h0e;
        mem[24] = 6'h05;
        mem[25] = 6'h3b;
        mem[26] = 6'h36;
        mem[27] = 6'h2d;
        mem[28] = 6'h3d;
        mem[29] = 6'h16;
        mem[30] = 6'h09;
        mem[31] = 6'h24;
        mem[32] = 6'h21;
        mem[33] = 6'h2c;
        mem[34] = 6'h2a;
        mem[35] = 6'h1a;
        mem[36] = 6'h30;
        mem[37] = 6'h0b;
        mem[38] = 6'h01;
        mem[39] = 6'h33;
        mem[40] = 6'h3f;
        mem[41] = 6'h39;
        mem[42] = 6'h23;
        mem[43] = 6'h15;
        mem[44] = 6'h02;
        mem[45] = 6'h20;
        mem[46] = 6'h3c;
        mem[47] = 6'h31;
        mem[48] = 6'h03;
        mem[49] = 6'h2b;
        mem[50] = 6'h1b;
        mem[51] = 6'h0c;
        mem[52] = 6'h3a;
        mem[53] = 6'h1f;
        mem[54] = 6'h0f;
        mem[55] = 6'h19;
        mem[56] = 6'h13;
        mem[57] = 6'h2e;
        mem[58] = 6'h11;
        mem[59] = 6'h0a;
        mem[60] = 6'h10;
        mem[61] = 6'h1c;
        mem[62] = 6'h04;
        mem[63] = 6'h22;
    end
endmodule

module encrypt_4sbox_large0(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h0d2;
        mem[1] = 10'h0f3;
        mem[2] = 10'h240;
        mem[3] = 10'h0d9;
        mem[4] = 10'h02d;
        mem[5] = 10'h33a;
        mem[6] = 10'h016;
        mem[7] = 10'h2af;
        mem[8] = 10'h0c8;
        mem[9] = 10'h224;
        mem[10] = 10'h3ec;
        mem[11] = 10'h14f;
        mem[12] = 10'h3d6;
        mem[13] = 10'h3ac;
        mem[14] = 10'h0a5;
        mem[15] = 10'h3ff;
        mem[16] = 10'h2a1;
        mem[17] = 10'h38d;
        mem[18] = 10'h3f2;
        mem[19] = 10'h2b8;
        mem[20] = 10'h3f9;
        mem[21] = 10'h243;
        mem[22] = 10'h30c;
        mem[23] = 10'h291;
        mem[24] = 10'h015;
        mem[25] = 10'h275;
        mem[26] = 10'h300;
        mem[27] = 10'h25a;
        mem[28] = 10'h221;
        mem[29] = 10'h389;
        mem[30] = 10'h13a;
        mem[31] = 10'h149;
        mem[32] = 10'h16c;
        mem[33] = 10'h2c3;
        mem[34] = 10'h117;
        mem[35] = 10'h305;
        mem[36] = 10'h020;
        mem[37] = 10'h14d;
        mem[38] = 10'h383;
        mem[39] = 10'h34b;
        mem[40] = 10'h381;
        mem[41] = 10'h25f;
        mem[42] = 10'h127;
        mem[43] = 10'h09f;
        mem[44] = 10'h292;
        mem[45] = 10'h027;
        mem[46] = 10'h29d;
        mem[47] = 10'h3c8;
        mem[48] = 10'h188;
        mem[49] = 10'h111;
        mem[50] = 10'h0f9;
        mem[51] = 10'h31d;
        mem[52] = 10'h023;
        mem[53] = 10'h355;
        mem[54] = 10'h2b0;
        mem[55] = 10'h33f;
        mem[56] = 10'h105;
        mem[57] = 10'h2de;
        mem[58] = 10'h191;
        mem[59] = 10'h1b5;
        mem[60] = 10'h27f;
        mem[61] = 10'h214;
        mem[62] = 10'h082;
        mem[63] = 10'h002;
        mem[64] = 10'h209;
        mem[65] = 10'h3ae;
        mem[66] = 10'h0e9;
        mem[67] = 10'h35e;
        mem[68] = 10'h1c2;
        mem[69] = 10'h177;
        mem[70] = 10'h047;
        mem[71] = 10'h0f7;
        mem[72] = 10'h03f;
        mem[73] = 10'h2bd;
        mem[74] = 10'h339;
        mem[75] = 10'h049;
        mem[76] = 10'h166;
        mem[77] = 10'h261;
        mem[78] = 10'h0b0;
        mem[79] = 10'h232;
        mem[80] = 10'h382;
        mem[81] = 10'h125;
        mem[82] = 10'h0db;
        mem[83] = 10'h000;
        mem[84] = 10'h070;
        mem[85] = 10'h3ce;
        mem[86] = 10'h343;
        mem[87] = 10'h1e6;
        mem[88] = 10'h35a;
        mem[89] = 10'h115;
        mem[90] = 10'h018;
        mem[91] = 10'h1bb;
        mem[92] = 10'h24e;
        mem[93] = 10'h38c;
        mem[94] = 10'h30b;
        mem[95] = 10'h201;
        mem[96] = 10'h1ed;
        mem[97] = 10'h306;
        mem[98] = 10'h233;
        mem[99] = 10'h137;
        mem[100] = 10'h290;
        mem[101] = 10'h3aa;
        mem[102] = 10'h187;
        mem[103] = 10'h212;
        mem[104] = 10'h37a;
        mem[105] = 10'h01e;
        mem[106] = 10'h0eb;
        mem[107] = 10'h1a8;
        mem[108] = 10'h3c5;
        mem[109] = 10'h13c;
        mem[110] = 10'h30a;
        mem[111] = 10'h039;
        mem[112] = 10'h2e8;
        mem[113] = 10'h0e6;
        mem[114] = 10'h3c2;
        mem[115] = 10'h3fa;
        mem[116] = 10'h124;
        mem[117] = 10'h025;
        mem[118] = 10'h078;
        mem[119] = 10'h29f;
        mem[120] = 10'h10f;
        mem[121] = 10'h0fe;
        mem[122] = 10'h349;
        mem[123] = 10'h2d4;
        mem[124] = 10'h0dc;
        mem[125] = 10'h150;
        mem[126] = 10'h216;
        mem[127] = 10'h277;
        mem[128] = 10'h2df;
        mem[129] = 10'h348;
        mem[130] = 10'h155;
        mem[131] = 10'h285;
        mem[132] = 10'h3de;
        mem[133] = 10'h3a9;
        mem[134] = 10'h3cb;
        mem[135] = 10'h1f3;
        mem[136] = 10'h378;
        mem[137] = 10'h2e3;
        mem[138] = 10'h1eb;
        mem[139] = 10'h06f;
        mem[140] = 10'h16b;
        mem[141] = 10'h2be;
        mem[142] = 10'h3be;
        mem[143] = 10'h2f8;
        mem[144] = 10'h07e;
        mem[145] = 10'h309;
        mem[146] = 10'h094;
        mem[147] = 10'h062;
        mem[148] = 10'h09a;
        mem[149] = 10'h058;
        mem[150] = 10'h2c2;
        mem[151] = 10'h1bc;
        mem[152] = 10'h0bd;
        mem[153] = 10'h0a0;
        mem[154] = 10'h04b;
        mem[155] = 10'h08c;
        mem[156] = 10'h20d;
        mem[157] = 10'h0a3;
        mem[158] = 10'h213;
        mem[159] = 10'h122;
        mem[160] = 10'h0ac;
        mem[161] = 10'h038;
        mem[162] = 10'h22a;
        mem[163] = 10'h283;
        mem[164] = 10'h251;
        mem[165] = 10'h2a7;
        mem[166] = 10'h026;
        mem[167] = 10'h079;
        mem[168] = 10'h0cc;
        mem[169] = 10'h156;
        mem[170] = 10'h02f;
        mem[171] = 10'h134;
        mem[172] = 10'h23d;
        mem[173] = 10'h1ee;
        mem[174] = 10'h1d3;
        mem[175] = 10'h100;
        mem[176] = 10'h21e;
        mem[177] = 10'h165;
        mem[178] = 10'h3e7;
        mem[179] = 10'h3db;
        mem[180] = 10'h225;
        mem[181] = 10'h199;
        mem[182] = 10'h266;
        mem[183] = 10'h318;
        mem[184] = 10'h351;
        mem[185] = 10'h257;
        mem[186] = 10'h3b5;
        mem[187] = 10'h271;
        mem[188] = 10'h121;
        mem[189] = 10'h29b;
        mem[190] = 10'h0a4;
        mem[191] = 10'h08f;
        mem[192] = 10'h3d7;
        mem[193] = 10'h106;
        mem[194] = 10'h15c;
        mem[195] = 10'h342;
        mem[196] = 10'h393;
        mem[197] = 10'h289;
        mem[198] = 10'h281;
        mem[199] = 10'h373;
        mem[200] = 10'h146;
        mem[201] = 10'h2f2;
        mem[202] = 10'h32e;
        mem[203] = 10'h1bd;
        mem[204] = 10'h31c;
        mem[205] = 10'h26c;
        mem[206] = 10'h264;
        mem[207] = 10'h0df;
        mem[208] = 10'h330;
        mem[209] = 10'h29a;
        mem[210] = 10'h024;
        mem[211] = 10'h314;
        mem[212] = 10'h129;
        mem[213] = 10'h05e;
        mem[214] = 10'h284;
        mem[215] = 10'h3ef;
        mem[216] = 10'h235;
        mem[217] = 10'h130;
        mem[218] = 10'h3bc;
        mem[219] = 10'h1cc;
        mem[220] = 10'h36a;
        mem[221] = 10'h04c;
        mem[222] = 10'h376;
        mem[223] = 10'h0ce;
        mem[224] = 10'h34a;
        mem[225] = 10'h21b;
        mem[226] = 10'h0c9;
        mem[227] = 10'h323;
        mem[228] = 10'h315;
        mem[229] = 10'h1a9;
        mem[230] = 10'h319;
        mem[231] = 10'h247;
        mem[232] = 10'h12f;
        mem[233] = 10'h0f6;
        mem[234] = 10'h11e;
        mem[235] = 10'h18c;
        mem[236] = 10'h1c1;
        mem[237] = 10'h006;
        mem[238] = 10'h13d;
        mem[239] = 10'h139;
        mem[240] = 10'h08e;
        mem[241] = 10'h365;
        mem[242] = 10'h26b;
        mem[243] = 10'h37f;
        mem[244] = 10'h2bc;
        mem[245] = 10'h089;
        mem[246] = 10'h0de;
        mem[247] = 10'h2b5;
        mem[248] = 10'h388;
        mem[249] = 10'h0d3;
        mem[250] = 10'h136;
        mem[251] = 10'h1b9;
        mem[252] = 10'h1e2;
        mem[253] = 10'h109;
        mem[254] = 10'h126;
        mem[255] = 10'h2ab;
        mem[256] = 10'h384;
        mem[257] = 10'h37b;
        mem[258] = 10'h157;
        mem[259] = 10'h3bf;
        mem[260] = 10'h19a;
        mem[261] = 10'h14b;
        mem[262] = 10'h068;
        mem[263] = 10'h0ba;
        mem[264] = 10'h1c4;
        mem[265] = 10'h1d7;
        mem[266] = 10'h238;
        mem[267] = 10'h14c;
        mem[268] = 10'h055;
        mem[269] = 10'h00a;
        mem[270] = 10'h10b;
        mem[271] = 10'h23e;
        mem[272] = 10'h043;
        mem[273] = 10'h24a;
        mem[274] = 10'h05f;
        mem[275] = 10'h2e0;
        mem[276] = 10'h311;
        mem[277] = 10'h084;
        mem[278] = 10'h175;
        mem[279] = 10'h06d;
        mem[280] = 10'h087;
        mem[281] = 10'h02a;
        mem[282] = 10'h242;
        mem[283] = 10'h3cd;
        mem[284] = 10'h37c;
        mem[285] = 10'h1cf;
        mem[286] = 10'h096;
        mem[287] = 10'h3d5;
        mem[288] = 10'h3fc;
        mem[289] = 10'h3e1;
        mem[290] = 10'h1b8;
        mem[291] = 10'h08a;
        mem[292] = 10'h215;
        mem[293] = 10'h190;
        mem[294] = 10'h3e5;
        mem[295] = 10'h138;
        mem[296] = 10'h3eb;
        mem[297] = 10'h2c1;
        mem[298] = 10'h2ac;
        mem[299] = 10'h1c3;
        mem[300] = 10'h218;
        mem[301] = 10'h3cf;
        mem[302] = 10'h0c0;
        mem[303] = 10'h06e;
        mem[304] = 10'h3e8;
        mem[305] = 10'h113;
        mem[306] = 10'h19c;
        mem[307] = 10'h317;
        mem[308] = 10'h202;
        mem[309] = 10'h052;
        mem[310] = 10'h09c;
        mem[311] = 10'h198;
        mem[312] = 10'h148;
        mem[313] = 10'h035;
        mem[314] = 10'h2ea;
        mem[315] = 10'h1fd;
        mem[316] = 10'h1aa;
        mem[317] = 10'h1c5;
        mem[318] = 10'h25d;
        mem[319] = 10'h010;
        mem[320] = 10'h13f;
        mem[321] = 10'h1ce;
        mem[322] = 10'h1be;
        mem[323] = 10'h30d;
        mem[324] = 10'h141;
        mem[325] = 10'h2eb;
        mem[326] = 10'h3b8;
        mem[327] = 10'h3af;
        mem[328] = 10'h0c1;
        mem[329] = 10'h11f;
        mem[330] = 10'h1d6;
        mem[331] = 10'h071;
        mem[332] = 10'h2b9;
        mem[333] = 10'h2d3;
        mem[334] = 10'h27c;
        mem[335] = 10'h1ec;
        mem[336] = 10'h0a2;
        mem[337] = 10'h178;
        mem[338] = 10'h0cd;
        mem[339] = 10'h120;
        mem[340] = 10'h02c;
        mem[341] = 10'h3d8;
        mem[342] = 10'h007;
        mem[343] = 10'h00d;
        mem[344] = 10'h0e4;
        mem[345] = 10'h0e1;
        mem[346] = 10'h227;
        mem[347] = 10'h3b3;
        mem[348] = 10'h142;
        mem[349] = 10'h174;
        mem[350] = 10'h2ee;
        mem[351] = 10'h143;
        mem[352] = 10'h2c7;
        mem[353] = 10'h12b;
        mem[354] = 10'h0af;
        mem[355] = 10'h0f0;
        mem[356] = 10'h1f8;
        mem[357] = 10'h0b7;
        mem[358] = 10'h046;
        mem[359] = 10'h255;
        mem[360] = 10'h107;
        mem[361] = 10'h0ca;
        mem[362] = 10'h164;
        mem[363] = 10'h152;
        mem[364] = 10'h075;
        mem[365] = 10'h3fe;
        mem[366] = 10'h23a;
        mem[367] = 10'h160;
        mem[368] = 10'h0cf;
        mem[369] = 10'h390;
        mem[370] = 10'h229;
        mem[371] = 10'h35b;
        mem[372] = 10'h01d;
        mem[373] = 10'h014;
        mem[374] = 10'h2ec;
        mem[375] = 10'h3ed;
        mem[376] = 10'h0d8;
        mem[377] = 10'h0c4;
        mem[378] = 10'h324;
        mem[379] = 10'h337;
        mem[380] = 10'h322;
        mem[381] = 10'h0f2;
        mem[382] = 10'h3b6;
        mem[383] = 10'h051;
        mem[384] = 10'h1dc;
        mem[385] = 10'h263;
        mem[386] = 10'h0d7;
        mem[387] = 10'h021;
        mem[388] = 10'h33b;
        mem[389] = 10'h0c2;
        mem[390] = 10'h1fc;
        mem[391] = 10'h02b;
        mem[392] = 10'h3f7;
        mem[393] = 10'h163;
        mem[394] = 10'h13b;
        mem[395] = 10'h3b9;
        mem[396] = 10'h1f1;
        mem[397] = 10'h3c0;
        mem[398] = 10'h326;
        mem[399] = 10'h350;
        mem[400] = 10'h207;
        mem[401] = 10'h293;
        mem[402] = 10'h2cd;
        mem[403] = 10'h282;
        mem[404] = 10'h369;
        mem[405] = 10'h2bf;
        mem[406] = 10'h3a8;
        mem[407] = 10'h1f9;
        mem[408] = 10'h108;
        mem[409] = 10'h162;
        mem[410] = 10'h17f;
        mem[411] = 10'h00c;
        mem[412] = 10'h245;
        mem[413] = 10'h1a7;
        mem[414] = 10'h06b;
        mem[415] = 10'h2da;
        mem[416] = 10'h1fb;
        mem[417] = 10'h222;
        mem[418] = 10'h2e4;
        mem[419] = 10'h280;
        mem[420] = 10'h045;
        mem[421] = 10'h3b1;
        mem[422] = 10'h39c;
        mem[423] = 10'h254;
        mem[424] = 10'h16d;
        mem[425] = 10'h03a;
        mem[426] = 10'h303;
        mem[427] = 10'h0b3;
        mem[428] = 10'h200;
        mem[429] = 10'h12c;
        mem[430] = 10'h09d;
        mem[431] = 10'h197;
        mem[432] = 10'h36c;
        mem[433] = 10'h0a6;
        mem[434] = 10'h04a;
        mem[435] = 10'h01a;
        mem[436] = 10'h29c;
        mem[437] = 10'h2b3;
        mem[438] = 10'h39a;
        mem[439] = 10'h27e;
        mem[440] = 10'h328;
        mem[441] = 10'h06c;
        mem[442] = 10'h308;
        mem[443] = 10'h0fc;
        mem[444] = 10'h325;
        mem[445] = 10'h25e;
        mem[446] = 10'h091;
        mem[447] = 10'h2fc;
        mem[448] = 10'h0c7;
        mem[449] = 10'h344;
        mem[450] = 10'h346;
        mem[451] = 10'h1e0;
        mem[452] = 10'h119;
        mem[453] = 10'h173;
        mem[454] = 10'h273;
        mem[455] = 10'h1df;
        mem[456] = 10'h042;
        mem[457] = 10'h1d8;
        mem[458] = 10'h16e;
        mem[459] = 10'h061;
        mem[460] = 10'h3bd;
        mem[461] = 10'h2f0;
        mem[462] = 10'h169;
        mem[463] = 10'h3b2;
        mem[464] = 10'h37e;
        mem[465] = 10'h09b;
        mem[466] = 10'h30e;
        mem[467] = 10'h0ff;
        mem[468] = 10'h2c8;
        mem[469] = 10'h272;
        mem[470] = 10'h26d;
        mem[471] = 10'h3e6;
        mem[472] = 10'h2fa;
        mem[473] = 10'h2d5;
        mem[474] = 10'h217;
        mem[475] = 10'h397;
        mem[476] = 10'h3dd;
        mem[477] = 10'h112;
        mem[478] = 10'h258;
        mem[479] = 10'h065;
        mem[480] = 10'h034;
        mem[481] = 10'h3f5;
        mem[482] = 10'h044;
        mem[483] = 10'h0b8;
        mem[484] = 10'h371;
        mem[485] = 10'h210;
        mem[486] = 10'h2dc;
        mem[487] = 10'h312;
        mem[488] = 10'h248;
        mem[489] = 10'h340;
        mem[490] = 10'h278;
        mem[491] = 10'h1ca;
        mem[492] = 10'h352;
        mem[493] = 10'h270;
        mem[494] = 10'h2c5;
        mem[495] = 10'h358;
        mem[496] = 10'h0f1;
        mem[497] = 10'h2d2;
        mem[498] = 10'h116;
        mem[499] = 10'h22d;
        mem[500] = 10'h181;
        mem[501] = 10'h063;
        mem[502] = 10'h056;
        mem[503] = 10'h377;
        mem[504] = 10'h1d9;
        mem[505] = 10'h360;
        mem[506] = 10'h183;
        mem[507] = 10'h20b;
        mem[508] = 10'h236;
        mem[509] = 10'h295;
        mem[510] = 10'h3b7;
        mem[511] = 10'h0ea;
        mem[512] = 10'h24d;
        mem[513] = 10'h3e3;
        mem[514] = 10'h004;
        mem[515] = 10'h3f4;
        mem[516] = 10'h170;
        mem[517] = 10'h32c;
        mem[518] = 10'h31e;
        mem[519] = 10'h21d;
        mem[520] = 10'h011;
        mem[521] = 10'h1dd;
        mem[522] = 10'h203;
        mem[523] = 10'h276;
        mem[524] = 10'h2f5;
        mem[525] = 10'h0e2;
        mem[526] = 10'h3fb;
        mem[527] = 10'h304;
        mem[528] = 10'h1da;
        mem[529] = 10'h118;
        mem[530] = 10'h101;
        mem[531] = 10'h39e;
        mem[532] = 10'h392;
        mem[533] = 10'h2d6;
        mem[534] = 10'h17a;
        mem[535] = 10'h2cf;
        mem[536] = 10'h060;
        mem[537] = 10'h20f;
        mem[538] = 10'h370;
        mem[539] = 10'h3c6;
        mem[540] = 10'h0c6;
        mem[541] = 10'h1cd;
        mem[542] = 10'h17b;
        mem[543] = 10'h083;
        mem[544] = 10'h1f4;
        mem[545] = 10'h18f;
        mem[546] = 10'h05d;
        mem[547] = 10'h25b;
        mem[548] = 10'h2d9;
        mem[549] = 10'h09e;
        mem[550] = 10'h246;
        mem[551] = 10'h32d;
        mem[552] = 10'h28b;
        mem[553] = 10'h15b;
        mem[554] = 10'h379;
        mem[555] = 10'h19f;
        mem[556] = 10'h03c;
        mem[557] = 10'h1d1;
        mem[558] = 10'h2dd;
        mem[559] = 10'h3f0;
        mem[560] = 10'h151;
        mem[561] = 10'h265;
        mem[562] = 10'h074;
        mem[563] = 10'h0b6;
        mem[564] = 10'h064;
        mem[565] = 10'h2e2;
        mem[566] = 10'h22e;
        mem[567] = 10'h0ee;
        mem[568] = 10'h24b;
        mem[569] = 10'h391;
        mem[570] = 10'h3d0;
        mem[571] = 10'h28c;
        mem[572] = 10'h103;
        mem[573] = 10'h208;
        mem[574] = 10'h17d;
        mem[575] = 10'h0ef;
        mem[576] = 10'h3dc;
        mem[577] = 10'h0f4;
        mem[578] = 10'h363;
        mem[579] = 10'h1ff;
        mem[580] = 10'h23f;
        mem[581] = 10'h3fd;
        mem[582] = 10'h1f5;
        mem[583] = 10'h037;
        mem[584] = 10'h294;
        mem[585] = 10'h2cb;
        mem[586] = 10'h1ef;
        mem[587] = 10'h1e9;
        mem[588] = 10'h2f4;
        mem[589] = 10'h3c1;
        mem[590] = 10'h2e1;
        mem[591] = 10'h19b;
        mem[592] = 10'h220;
        mem[593] = 10'h25c;
        mem[594] = 10'h0c3;
        mem[595] = 10'h00f;
        mem[596] = 10'h06a;
        mem[597] = 10'h3e4;
        mem[598] = 10'h158;
        mem[599] = 10'h234;
        mem[600] = 10'h356;
        mem[601] = 10'h036;
        mem[602] = 10'h01c;
        mem[603] = 10'h3d2;
        mem[604] = 10'h0e0;
        mem[605] = 10'h3da;
        mem[606] = 10'h335;
        mem[607] = 10'h3ca;
        mem[608] = 10'h171;
        mem[609] = 10'h34d;
        mem[610] = 10'h239;
        mem[611] = 10'h080;
        mem[612] = 10'h19d;
        mem[613] = 10'h3d4;
        mem[614] = 10'h0b4;
        mem[615] = 10'h3d3;
        mem[616] = 10'h147;
        mem[617] = 10'h2e7;
        mem[618] = 10'h35c;
        mem[619] = 10'h040;
        mem[620] = 10'h005;
        mem[621] = 10'h2f9;
        mem[622] = 10'h0be;
        mem[623] = 10'h1f7;
        mem[624] = 10'h0d6;
        mem[625] = 10'h00e;
        mem[626] = 10'h0fd;
        mem[627] = 10'h1db;
        mem[628] = 10'h3f1;
        mem[629] = 10'h2ed;
        mem[630] = 10'h067;
        mem[631] = 10'h0bf;
        mem[632] = 10'h38a;
        mem[633] = 10'h29e;
        mem[634] = 10'h04d;
        mem[635] = 10'h0b5;
        mem[636] = 10'h001;
        mem[637] = 10'h069;
        mem[638] = 10'h172;
        mem[639] = 10'h396;
        mem[640] = 10'h1b2;
        mem[641] = 10'h05b;
        mem[642] = 10'h2e5;
        mem[643] = 10'h185;
        mem[644] = 10'h031;
        mem[645] = 10'h0aa;
        mem[646] = 10'h2ff;
        mem[647] = 10'h299;
        mem[648] = 10'h189;
        mem[649] = 10'h18a;
        mem[650] = 10'h250;
        mem[651] = 10'h1f6;
        mem[652] = 10'h38b;
        mem[653] = 10'h0fb;
        mem[654] = 10'h050;
        mem[655] = 10'h3c9;
        mem[656] = 10'h3a1;
        mem[657] = 10'h003;
        mem[658] = 10'h316;
        mem[659] = 10'h1f0;
        mem[660] = 10'h361;
        mem[661] = 10'h05a;
        mem[662] = 10'h18e;
        mem[663] = 10'h353;
        mem[664] = 10'h15e;
        mem[665] = 10'h073;
        mem[666] = 10'h1a1;
        mem[667] = 10'h3b4;
        mem[668] = 10'h08d;
        mem[669] = 10'h32a;
        mem[670] = 10'h3a0;
        mem[671] = 10'h2b6;
        mem[672] = 10'h2c4;
        mem[673] = 10'h36f;
        mem[674] = 10'h15f;
        mem[675] = 10'h3e9;
        mem[676] = 10'h16f;
        mem[677] = 10'h338;
        mem[678] = 10'h387;
        mem[679] = 10'h321;
        mem[680] = 10'h008;
        mem[681] = 10'h2e9;
        mem[682] = 10'h03e;
        mem[683] = 10'h2bb;
        mem[684] = 10'h28f;
        mem[685] = 10'h367;
        mem[686] = 10'h095;
        mem[687] = 10'h366;
        mem[688] = 10'h2ba;
        mem[689] = 10'h34c;
        mem[690] = 10'h022;
        mem[691] = 10'h341;
        mem[692] = 10'h133;
        mem[693] = 10'h098;
        mem[694] = 10'h07f;
        mem[695] = 10'h18d;
        mem[696] = 10'h12a;
        mem[697] = 10'h24f;
        mem[698] = 10'h140;
        mem[699] = 10'h092;
        mem[700] = 10'h33c;
        mem[701] = 10'h0bb;
        mem[702] = 10'h0ab;
        mem[703] = 10'h226;
        mem[704] = 10'h15d;
        mem[705] = 10'h161;
        mem[706] = 10'h3ba;
        mem[707] = 10'h1c0;
        mem[708] = 10'h35d;
        mem[709] = 10'h132;
        mem[710] = 10'h1b4;
        mem[711] = 10'h07b;
        mem[712] = 10'h11a;
        mem[713] = 10'h07a;
        mem[714] = 10'h17c;
        mem[715] = 10'h10a;
        mem[716] = 10'h21c;
        mem[717] = 10'h347;
        mem[718] = 10'h1ab;
        mem[719] = 10'h2a0;
        mem[720] = 10'h10e;
        mem[721] = 10'h36d;
        mem[722] = 10'h3f3;
        mem[723] = 10'h231;
        mem[724] = 10'h374;
        mem[725] = 10'h27d;
        mem[726] = 10'h0ad;
        mem[727] = 10'h0a9;
        mem[728] = 10'h20a;
        mem[729] = 10'h08b;
        mem[730] = 10'h375;
        mem[731] = 10'h176;
        mem[732] = 10'h12e;
        mem[733] = 10'h1d5;
        mem[734] = 10'h10d;
        mem[735] = 10'h20c;
        mem[736] = 10'h354;
        mem[737] = 10'h380;
        mem[738] = 10'h0d5;
        mem[739] = 10'h252;
        mem[740] = 10'h0a7;
        mem[741] = 10'h1a5;
        mem[742] = 10'h260;
        mem[743] = 10'h009;
        mem[744] = 10'h39f;
        mem[745] = 10'h1fa;
        mem[746] = 10'h088;
        mem[747] = 10'h205;
        mem[748] = 10'h3a6;
        mem[749] = 10'h3ea;
        mem[750] = 10'h334;
        mem[751] = 10'h394;
        mem[752] = 10'h38e;
        mem[753] = 10'h241;
        mem[754] = 10'h3c3;
        mem[755] = 10'h07c;
        mem[756] = 10'h26e;
        mem[757] = 10'h2ae;
        mem[758] = 10'h153;
        mem[759] = 10'h286;
        mem[760] = 10'h287;
        mem[761] = 10'h012;
        mem[762] = 10'h1b1;
        mem[763] = 10'h1de;
        mem[764] = 10'h1ac;
        mem[765] = 10'h0bc;
        mem[766] = 10'h192;
        mem[767] = 10'h0d1;
        mem[768] = 10'h3ee;
        mem[769] = 10'h013;
        mem[770] = 10'h3bb;
        mem[771] = 10'h2d0;
        mem[772] = 10'h36e;
        mem[773] = 10'h336;
        mem[774] = 10'h2d7;
        mem[775] = 10'h357;
        mem[776] = 10'h2db;
        mem[777] = 10'h307;
        mem[778] = 10'h029;
        mem[779] = 10'h2a8;
        mem[780] = 10'h2aa;
        mem[781] = 10'h345;
        mem[782] = 10'h085;
        mem[783] = 10'h329;
        mem[784] = 10'h0a1;
        mem[785] = 10'h3f8;
        mem[786] = 10'h22f;
        mem[787] = 10'h1a4;
        mem[788] = 10'h194;
        mem[789] = 10'h2b4;
        mem[790] = 10'h033;
        mem[791] = 10'h1f2;
        mem[792] = 10'h39d;
        mem[793] = 10'h14e;
        mem[794] = 10'h1e5;
        mem[795] = 10'h2a9;
        mem[796] = 10'h288;
        mem[797] = 10'h0f8;
        mem[798] = 10'h206;
        mem[799] = 10'h131;
        mem[800] = 10'h2a3;
        mem[801] = 10'h368;
        mem[802] = 10'h2d1;
        mem[803] = 10'h02e;
        mem[804] = 10'h1a6;
        mem[805] = 10'h07d;
        mem[806] = 10'h03b;
        mem[807] = 10'h12d;
        mem[808] = 10'h3ab;
        mem[809] = 10'h230;
        mem[810] = 10'h1a3;
        mem[811] = 10'h36b;
        mem[812] = 10'h223;
        mem[813] = 10'h3df;
        mem[814] = 10'h0e5;
        mem[815] = 10'h0d4;
        mem[816] = 10'h144;
        mem[817] = 10'h196;
        mem[818] = 10'h301;
        mem[819] = 10'h11d;
        mem[820] = 10'h1bf;
        mem[821] = 10'h320;
        mem[822] = 10'h2b2;
        mem[823] = 10'h072;
        mem[824] = 10'h0da;
        mem[825] = 10'h267;
        mem[826] = 10'h2fd;
        mem[827] = 10'h26a;
        mem[828] = 10'h385;
        mem[829] = 10'h32f;
        mem[830] = 10'h3e2;
        mem[831] = 10'h04e;
        mem[832] = 10'h33e;
        mem[833] = 10'h1e1;
        mem[834] = 10'h359;
        mem[835] = 10'h364;
        mem[836] = 10'h398;
        mem[837] = 10'h2a6;
        mem[838] = 10'h066;
        mem[839] = 10'h2ce;
        mem[840] = 10'h3b0;
        mem[841] = 10'h00b;
        mem[842] = 10'h1cb;
        mem[843] = 10'h3c4;
        mem[844] = 10'h31a;
        mem[845] = 10'h2ef;
        mem[846] = 10'h253;
        mem[847] = 10'h04f;
        mem[848] = 10'h01f;
        mem[849] = 10'h27b;
        mem[850] = 10'h28d;
        mem[851] = 10'h2d8;
        mem[852] = 10'h1fe;
        mem[853] = 10'h053;
        mem[854] = 10'h269;
        mem[855] = 10'h05c;
        mem[856] = 10'h1b7;
        mem[857] = 10'h296;
        mem[858] = 10'h34f;
        mem[859] = 10'h32b;
        mem[860] = 10'h26f;
        mem[861] = 10'h099;
        mem[862] = 10'h1d2;
        mem[863] = 10'h1b3;
        mem[864] = 10'h102;
        mem[865] = 10'h017;
        mem[866] = 10'h11c;
        mem[867] = 10'h332;
        mem[868] = 10'h0e8;
        mem[869] = 10'h159;
        mem[870] = 10'h3d9;
        mem[871] = 10'h298;
        mem[872] = 10'h195;
        mem[873] = 10'h081;
        mem[874] = 10'h37d;
        mem[875] = 10'h327;
        mem[876] = 10'h3c7;
        mem[877] = 10'h168;
        mem[878] = 10'h2c9;
        mem[879] = 10'h0fa;
        mem[880] = 10'h1e7;
        mem[881] = 10'h2e6;
        mem[882] = 10'h2a2;
        mem[883] = 10'h2fe;
        mem[884] = 10'h33d;
        mem[885] = 10'h1ea;
        mem[886] = 10'h39b;
        mem[887] = 10'h11b;
        mem[888] = 10'h34e;
        mem[889] = 10'h0ae;
        mem[890] = 10'h1c8;
        mem[891] = 10'h048;
        mem[892] = 10'h268;
        mem[893] = 10'h154;
        mem[894] = 10'h0e7;
        mem[895] = 10'h24c;
        mem[896] = 10'h31b;
        mem[897] = 10'h1b0;
        mem[898] = 10'h1c6;
        mem[899] = 10'h13e;
        mem[900] = 10'h0a8;
        mem[901] = 10'h21a;
        mem[902] = 10'h193;
        mem[903] = 10'h2cc;
        mem[904] = 10'h2a4;
        mem[905] = 10'h1c9;
        mem[906] = 10'h395;
        mem[907] = 10'h362;
        mem[908] = 10'h059;
        mem[909] = 10'h3a3;
        mem[910] = 10'h032;
        mem[911] = 10'h1b6;
        mem[912] = 10'h3f6;
        mem[913] = 10'h2f3;
        mem[914] = 10'h054;
        mem[915] = 10'h3cc;
        mem[916] = 10'h0b9;
        mem[917] = 10'h2c6;
        mem[918] = 10'h0f5;
        mem[919] = 10'h01b;
        mem[920] = 10'h128;
        mem[921] = 10'h21f;
        mem[922] = 10'h262;
        mem[923] = 10'h228;
        mem[924] = 10'h2f6;
        mem[925] = 10'h077;
        mem[926] = 10'h0c5;
        mem[927] = 10'h3ad;
        mem[928] = 10'h03d;
        mem[929] = 10'h3a2;
        mem[930] = 10'h1af;
        mem[931] = 10'h167;
        mem[932] = 10'h123;
        mem[933] = 10'h22c;
        mem[934] = 10'h086;
        mem[935] = 10'h1a0;
        mem[936] = 10'h22b;
        mem[937] = 10'h3e0;
        mem[938] = 10'h135;
        mem[939] = 10'h23c;
        mem[940] = 10'h3a5;
        mem[941] = 10'h2a5;
        mem[942] = 10'h219;
        mem[943] = 10'h1e4;
        mem[944] = 10'h331;
        mem[945] = 10'h399;
        mem[946] = 10'h057;
        mem[947] = 10'h302;
        mem[948] = 10'h249;
        mem[949] = 10'h10c;
        mem[950] = 10'h0cb;
        mem[951] = 10'h279;
        mem[952] = 10'h2ca;
        mem[953] = 10'h27a;
        mem[954] = 10'h310;
        mem[955] = 10'h19e;
        mem[956] = 10'h20e;
        mem[957] = 10'h2b7;
        mem[958] = 10'h179;
        mem[959] = 10'h041;
        mem[960] = 10'h0b2;
        mem[961] = 10'h35f;
        mem[962] = 10'h30f;
        mem[963] = 10'h333;
        mem[964] = 10'h184;
        mem[965] = 10'h180;
        mem[966] = 10'h1c7;
        mem[967] = 10'h2fb;
        mem[968] = 10'h2f1;
        mem[969] = 10'h076;
        mem[970] = 10'h0b1;
        mem[971] = 10'h244;
        mem[972] = 10'h1ba;
        mem[973] = 10'h1ae;
        mem[974] = 10'h097;
        mem[975] = 10'h38f;
        mem[976] = 10'h1d0;
        mem[977] = 10'h0d0;
        mem[978] = 10'h2ad;
        mem[979] = 10'h104;
        mem[980] = 10'h0ec;
        mem[981] = 10'h090;
        mem[982] = 10'h204;
        mem[983] = 10'h16a;
        mem[984] = 10'h237;
        mem[985] = 10'h3a7;
        mem[986] = 10'h17e;
        mem[987] = 10'h0e3;
        mem[988] = 10'h31f;
        mem[989] = 10'h28e;
        mem[990] = 10'h2f7;
        mem[991] = 10'h1d4;
        mem[992] = 10'h3d1;
        mem[993] = 10'h386;
        mem[994] = 10'h145;
        mem[995] = 10'h313;
        mem[996] = 10'h182;
        mem[997] = 10'h28a;
        mem[998] = 10'h1ad;
        mem[999] = 10'h259;
        mem[1000] = 10'h211;
        mem[1001] = 10'h093;
        mem[1002] = 10'h372;
        mem[1003] = 10'h0dd;
        mem[1004] = 10'h019;
        mem[1005] = 10'h14a;
        mem[1006] = 10'h1a2;
        mem[1007] = 10'h274;
        mem[1008] = 10'h18b;
        mem[1009] = 10'h030;
        mem[1010] = 10'h2b1;
        mem[1011] = 10'h1e8;
        mem[1012] = 10'h297;
        mem[1013] = 10'h256;
        mem[1014] = 10'h2c0;
        mem[1015] = 10'h23b;
        mem[1016] = 10'h15a;
        mem[1017] = 10'h1e3;
        mem[1018] = 10'h0ed;
        mem[1019] = 10'h114;
        mem[1020] = 10'h3a4;
        mem[1021] = 10'h110;
        mem[1022] = 10'h028;
        mem[1023] = 10'h186;
    end
endmodule

module encrypt_4sbox_large1(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h237;
        mem[1] = 10'h256;
        mem[2] = 10'h14e;
        mem[3] = 10'h166;
        mem[4] = 10'h048;
        mem[5] = 10'h1eb;
        mem[6] = 10'h240;
        mem[7] = 10'h2bd;
        mem[8] = 10'h129;
        mem[9] = 10'h2fa;
        mem[10] = 10'h38d;
        mem[11] = 10'h016;
        mem[12] = 10'h1da;
        mem[13] = 10'h2c9;
        mem[14] = 10'h0dd;
        mem[15] = 10'h2f7;
        mem[16] = 10'h1a0;
        mem[17] = 10'h3a0;
        mem[18] = 10'h3c1;
        mem[19] = 10'h0e9;
        mem[20] = 10'h1aa;
        mem[21] = 10'h394;
        mem[22] = 10'h1af;
        mem[23] = 10'h378;
        mem[24] = 10'h021;
        mem[25] = 10'h1d5;
        mem[26] = 10'h299;
        mem[27] = 10'h23c;
        mem[28] = 10'h23b;
        mem[29] = 10'h093;
        mem[30] = 10'h249;
        mem[31] = 10'h211;
        mem[32] = 10'h175;
        mem[33] = 10'h06e;
        mem[34] = 10'h123;
        mem[35] = 10'h24f;
        mem[36] = 10'h0cd;
        mem[37] = 10'h253;
        mem[38] = 10'h1ff;
        mem[39] = 10'h050;
        mem[40] = 10'h32d;
        mem[41] = 10'h00e;
        mem[42] = 10'h34d;
        mem[43] = 10'h05e;
        mem[44] = 10'h280;
        mem[45] = 10'h099;
        mem[46] = 10'h3c5;
        mem[47] = 10'h372;
        mem[48] = 10'h221;
        mem[49] = 10'h18e;
        mem[50] = 10'h2c7;
        mem[51] = 10'h3f1;
        mem[52] = 10'h008;
        mem[53] = 10'h2e9;
        mem[54] = 10'h01c;
        mem[55] = 10'h0bb;
        mem[56] = 10'h122;
        mem[57] = 10'h27f;
        mem[58] = 10'h132;
        mem[59] = 10'h1bc;
        mem[60] = 10'h0f6;
        mem[61] = 10'h33e;
        mem[62] = 10'h03d;
        mem[63] = 10'h374;
        mem[64] = 10'h2c4;
        mem[65] = 10'h3f0;
        mem[66] = 10'h164;
        mem[67] = 10'h2aa;
        mem[68] = 10'h281;
        mem[69] = 10'h07b;
        mem[70] = 10'h2f3;
        mem[71] = 10'h201;
        mem[72] = 10'h13a;
        mem[73] = 10'h2ae;
        mem[74] = 10'h0cc;
        mem[75] = 10'h02e;
        mem[76] = 10'h03c;
        mem[77] = 10'h1c9;
        mem[78] = 10'h2ce;
        mem[79] = 10'h0d1;
        mem[80] = 10'h30e;
        mem[81] = 10'h30d;
        mem[82] = 10'h058;
        mem[83] = 10'h0ed;
        mem[84] = 10'h335;
        mem[85] = 10'h257;
        mem[86] = 10'h3ab;
        mem[87] = 10'h0b3;
        mem[88] = 10'h112;
        mem[89] = 10'h3a2;
        mem[90] = 10'h31a;
        mem[91] = 10'h250;
        mem[92] = 10'h07d;
        mem[93] = 10'h29d;
        mem[94] = 10'h283;
        mem[95] = 10'h26c;
        mem[96] = 10'h219;
        mem[97] = 10'h3ac;
        mem[98] = 10'h37c;
        mem[99] = 10'h1b8;
        mem[100] = 10'h0dc;
        mem[101] = 10'h09b;
        mem[102] = 10'h37d;
        mem[103] = 10'h320;
        mem[104] = 10'h1a4;
        mem[105] = 10'h054;
        mem[106] = 10'h172;
        mem[107] = 10'h239;
        mem[108] = 10'h32e;
        mem[109] = 10'h1dd;
        mem[110] = 10'h326;
        mem[111] = 10'h210;
        mem[112] = 10'h03f;
        mem[113] = 10'h020;
        mem[114] = 10'h12f;
        mem[115] = 10'h0c4;
        mem[116] = 10'h080;
        mem[117] = 10'h3d6;
        mem[118] = 10'h024;
        mem[119] = 10'h2b3;
        mem[120] = 10'h365;
        mem[121] = 10'h139;
        mem[122] = 10'h03b;
        mem[123] = 10'h332;
        mem[124] = 10'h25c;
        mem[125] = 10'h35f;
        mem[126] = 10'h08e;
        mem[127] = 10'h011;
        mem[128] = 10'h2da;
        mem[129] = 10'h21c;
        mem[130] = 10'h1ae;
        mem[131] = 10'h247;
        mem[132] = 10'h2f9;
        mem[133] = 10'h2ad;
        mem[134] = 10'h387;
        mem[135] = 10'h1e7;
        mem[136] = 10'h346;
        mem[137] = 10'h012;
        mem[138] = 10'h2d0;
        mem[139] = 10'h342;
        mem[140] = 10'h36d;
        mem[141] = 10'h109;
        mem[142] = 10'h026;
        mem[143] = 10'h1f7;
        mem[144] = 10'h3e3;
        mem[145] = 10'h32a;
        mem[146] = 10'h3ba;
        mem[147] = 10'h0e1;
        mem[148] = 10'h176;
        mem[149] = 10'h3c4;
        mem[150] = 10'h0a6;
        mem[151] = 10'h1ee;
        mem[152] = 10'h186;
        mem[153] = 10'h00f;
        mem[154] = 10'h0f2;
        mem[155] = 10'h2ab;
        mem[156] = 10'h1fd;
        mem[157] = 10'h3e7;
        mem[158] = 10'h265;
        mem[159] = 10'h0ba;
        mem[160] = 10'h2a0;
        mem[161] = 10'h0eb;
        mem[162] = 10'h3cb;
        mem[163] = 10'h347;
        mem[164] = 10'h2e5;
        mem[165] = 10'h2cd;
        mem[166] = 10'h114;
        mem[167] = 10'h06f;
        mem[168] = 10'h036;
        mem[169] = 10'h10b;
        mem[170] = 10'h027;
        mem[171] = 10'h355;
        mem[172] = 10'h06b;
        mem[173] = 10'h11c;
        mem[174] = 10'h0f1;
        mem[175] = 10'h3c2;
        mem[176] = 10'h354;
        mem[177] = 10'h08b;
        mem[178] = 10'h17d;
        mem[179] = 10'h052;
        mem[180] = 10'h327;
        mem[181] = 10'h3d0;
        mem[182] = 10'h3db;
        mem[183] = 10'h18f;
        mem[184] = 10'h137;
        mem[185] = 10'h3fd;
        mem[186] = 10'h33a;
        mem[187] = 10'h1c7;
        mem[188] = 10'h1b4;
        mem[189] = 10'h125;
        mem[190] = 10'h2bc;
        mem[191] = 10'h343;
        mem[192] = 10'h0e2;
        mem[193] = 10'h15c;
        mem[194] = 10'h2be;
        mem[195] = 10'h0e6;
        mem[196] = 10'h15d;
        mem[197] = 10'h3cc;
        mem[198] = 10'h046;
        mem[199] = 10'h14b;
        mem[200] = 10'h205;
        mem[201] = 10'h2e1;
        mem[202] = 10'h1a6;
        mem[203] = 10'h315;
        mem[204] = 10'h1bf;
        mem[205] = 10'h0de;
        mem[206] = 10'h13b;
        mem[207] = 10'h1db;
        mem[208] = 10'h076;
        mem[209] = 10'h1c4;
        mem[210] = 10'h05c;
        mem[211] = 10'h282;
        mem[212] = 10'h0e8;
        mem[213] = 10'h2d8;
        mem[214] = 10'h0c9;
        mem[215] = 10'h3a1;
        mem[216] = 10'h185;
        mem[217] = 10'h1f0;
        mem[218] = 10'h2b7;
        mem[219] = 10'h073;
        mem[220] = 10'h35a;
        mem[221] = 10'h392;
        mem[222] = 10'h017;
        mem[223] = 10'h3be;
        mem[224] = 10'h3e2;
        mem[225] = 10'h1b5;
        mem[226] = 10'h2fc;
        mem[227] = 10'h36c;
        mem[228] = 10'h1b7;
        mem[229] = 10'h0c3;
        mem[230] = 10'h0d4;
        mem[231] = 10'h119;
        mem[232] = 10'h23e;
        mem[233] = 10'h015;
        mem[234] = 10'h2ee;
        mem[235] = 10'h0a2;
        mem[236] = 10'h2a8;
        mem[237] = 10'h26a;
        mem[238] = 10'h31e;
        mem[239] = 10'h095;
        mem[240] = 10'h181;
        mem[241] = 10'h2c5;
        mem[242] = 10'h07c;
        mem[243] = 10'h1a2;
        mem[244] = 10'h3dd;
        mem[245] = 10'h11a;
        mem[246] = 10'h0ea;
        mem[247] = 10'h005;
        mem[248] = 10'h36e;
        mem[249] = 10'h3da;
        mem[250] = 10'h255;
        mem[251] = 10'h041;
        mem[252] = 10'h2c0;
        mem[253] = 10'h149;
        mem[254] = 10'h1ca;
        mem[255] = 10'h353;
        mem[256] = 10'h2fe;
        mem[257] = 10'h0fe;
        mem[258] = 10'h1e4;
        mem[259] = 10'h1f8;
        mem[260] = 10'h31b;
        mem[261] = 10'h328;
        mem[262] = 10'h3bd;
        mem[263] = 10'h26b;
        mem[264] = 10'h3ea;
        mem[265] = 10'h316;
        mem[266] = 10'h23f;
        mem[267] = 10'h13c;
        mem[268] = 10'h07f;
        mem[269] = 10'h167;
        mem[270] = 10'h01b;
        mem[271] = 10'h307;
        mem[272] = 10'h1c2;
        mem[273] = 10'h0ae;
        mem[274] = 10'h27a;
        mem[275] = 10'h01f;
        mem[276] = 10'h1c8;
        mem[277] = 10'h2e4;
        mem[278] = 10'h13f;
        mem[279] = 10'h1d9;
        mem[280] = 10'h1ad;
        mem[281] = 10'h14f;
        mem[282] = 10'h0a7;
        mem[283] = 10'h33c;
        mem[284] = 10'h269;
        mem[285] = 10'h359;
        mem[286] = 10'h3d8;
        mem[287] = 10'h177;
        mem[288] = 10'h27e;
        mem[289] = 10'h364;
        mem[290] = 10'h1d7;
        mem[291] = 10'h01a;
        mem[292] = 10'h169;
        mem[293] = 10'h1a1;
        mem[294] = 10'h3c8;
        mem[295] = 10'h104;
        mem[296] = 10'h31c;
        mem[297] = 10'h04a;
        mem[298] = 10'h1cc;
        mem[299] = 10'h264;
        mem[300] = 10'h385;
        mem[301] = 10'h3b8;
        mem[302] = 10'h206;
        mem[303] = 10'h2f0;
        mem[304] = 10'h05b;
        mem[305] = 10'h218;
        mem[306] = 10'h187;
        mem[307] = 10'h0a3;
        mem[308] = 10'h3b2;
        mem[309] = 10'h3df;
        mem[310] = 10'h2a9;
        mem[311] = 10'h375;
        mem[312] = 10'h2ac;
        mem[313] = 10'h089;
        mem[314] = 10'h154;
        mem[315] = 10'h305;
        mem[316] = 10'h2e8;
        mem[317] = 10'h106;
        mem[318] = 10'h226;
        mem[319] = 10'h0c5;
        mem[320] = 10'h0ad;
        mem[321] = 10'h0c7;
        mem[322] = 10'h32c;
        mem[323] = 10'h0f0;
        mem[324] = 10'h2cb;
        mem[325] = 10'h303;
        mem[326] = 10'h35e;
        mem[327] = 10'h147;
        mem[328] = 10'h142;
        mem[329] = 10'h00a;
        mem[330] = 10'h3aa;
        mem[331] = 10'h2d3;
        mem[332] = 10'h0f3;
        mem[333] = 10'h18a;
        mem[334] = 10'h088;
        mem[335] = 10'h145;
        mem[336] = 10'h146;
        mem[337] = 10'h379;
        mem[338] = 10'h1ce;
        mem[339] = 10'h0b0;
        mem[340] = 10'h037;
        mem[341] = 10'h20d;
        mem[342] = 10'h203;
        mem[343] = 10'h17b;
        mem[344] = 10'h34e;
        mem[345] = 10'h00c;
        mem[346] = 10'h3e9;
        mem[347] = 10'h297;
        mem[348] = 10'h06d;
        mem[349] = 10'h2dd;
        mem[350] = 10'h28f;
        mem[351] = 10'h3ee;
        mem[352] = 10'h0f7;
        mem[353] = 10'h28a;
        mem[354] = 10'h25d;
        mem[355] = 10'h200;
        mem[356] = 10'h258;
        mem[357] = 10'h117;
        mem[358] = 10'h0f9;
        mem[359] = 10'h348;
        mem[360] = 10'h1de;
        mem[361] = 10'h049;
        mem[362] = 10'h22a;
        mem[363] = 10'h06c;
        mem[364] = 10'h213;
        mem[365] = 10'h3ad;
        mem[366] = 10'h216;
        mem[367] = 10'h196;
        mem[368] = 10'h276;
        mem[369] = 10'h2ba;
        mem[370] = 10'h0ce;
        mem[371] = 10'h014;
        mem[372] = 10'h301;
        mem[373] = 10'h031;
        mem[374] = 10'h032;
        mem[375] = 10'h22e;
        mem[376] = 10'h304;
        mem[377] = 10'h2d4;
        mem[378] = 10'h1a3;
        mem[379] = 10'h1fc;
        mem[380] = 10'h204;
        mem[381] = 10'h0d8;
        mem[382] = 10'h0d7;
        mem[383] = 10'h0e5;
        mem[384] = 10'h3b0;
        mem[385] = 10'h022;
        mem[386] = 10'h34c;
        mem[387] = 10'h383;
        mem[388] = 10'h1d1;
        mem[389] = 10'h370;
        mem[390] = 10'h143;
        mem[391] = 10'h3b4;
        mem[392] = 10'h092;
        mem[393] = 10'h1c5;
        mem[394] = 10'h231;
        mem[395] = 10'h292;
        mem[396] = 10'h188;
        mem[397] = 10'h3ec;
        mem[398] = 10'h386;
        mem[399] = 10'h3e5;
        mem[400] = 10'h01e;
        mem[401] = 10'h0e3;
        mem[402] = 10'h056;
        mem[403] = 10'h314;
        mem[404] = 10'h289;
        mem[405] = 10'h2c2;
        mem[406] = 10'h0d3;
        mem[407] = 10'h215;
        mem[408] = 10'h08a;
        mem[409] = 10'h11b;
        mem[410] = 10'h3d3;
        mem[411] = 10'h006;
        mem[412] = 10'h338;
        mem[413] = 10'h111;
        mem[414] = 10'h38b;
        mem[415] = 10'h09e;
        mem[416] = 10'h3e0;
        mem[417] = 10'h1c3;
        mem[418] = 10'h0f4;
        mem[419] = 10'h3e4;
        mem[420] = 10'h2b1;
        mem[421] = 10'h300;
        mem[422] = 10'h3fb;
        mem[423] = 10'h16a;
        mem[424] = 10'h018;
        mem[425] = 10'h37b;
        mem[426] = 10'h2a1;
        mem[427] = 10'h333;
        mem[428] = 10'h20b;
        mem[429] = 10'h057;
        mem[430] = 10'h086;
        mem[431] = 10'h2b4;
        mem[432] = 10'h3d1;
        mem[433] = 10'h2ca;
        mem[434] = 10'h0d2;
        mem[435] = 10'h0fa;
        mem[436] = 10'h34f;
        mem[437] = 10'h389;
        mem[438] = 10'h2ff;
        mem[439] = 10'h2c6;
        mem[440] = 10'h3fc;
        mem[441] = 10'h3ff;
        mem[442] = 10'h0fd;
        mem[443] = 10'h08f;
        mem[444] = 10'h1f5;
        mem[445] = 10'h159;
        mem[446] = 10'h232;
        mem[447] = 10'h0e0;
        mem[448] = 10'h199;
        mem[449] = 10'h2d7;
        mem[450] = 10'h39b;
        mem[451] = 10'h11d;
        mem[452] = 10'h242;
        mem[453] = 10'h3f5;
        mem[454] = 10'h29b;
        mem[455] = 10'h1f9;
        mem[456] = 10'h295;
        mem[457] = 10'h182;
        mem[458] = 10'h296;
        mem[459] = 10'h1cb;
        mem[460] = 10'h115;
        mem[461] = 10'h3d2;
        mem[462] = 10'h2b2;
        mem[463] = 10'h083;
        mem[464] = 10'h152;
        mem[465] = 10'h310;
        mem[466] = 10'h1a7;
        mem[467] = 10'h2c1;
        mem[468] = 10'h04b;
        mem[469] = 10'h28e;
        mem[470] = 10'h1a9;
        mem[471] = 10'h357;
        mem[472] = 10'h312;
        mem[473] = 10'h278;
        mem[474] = 10'h368;
        mem[475] = 10'h33f;
        mem[476] = 10'h0d0;
        mem[477] = 10'h1c0;
        mem[478] = 10'h286;
        mem[479] = 10'h3bf;
        mem[480] = 10'h2f4;
        mem[481] = 10'h329;
        mem[482] = 10'h2a6;
        mem[483] = 10'h0d5;
        mem[484] = 10'h11f;
        mem[485] = 10'h04f;
        mem[486] = 10'h17f;
        mem[487] = 10'h0e4;
        mem[488] = 10'h195;
        mem[489] = 10'h0f8;
        mem[490] = 10'h191;
        mem[491] = 10'h15f;
        mem[492] = 10'h127;
        mem[493] = 10'h261;
        mem[494] = 10'h271;
        mem[495] = 10'h352;
        mem[496] = 10'h044;
        mem[497] = 10'h192;
        mem[498] = 10'h071;
        mem[499] = 10'h294;
        mem[500] = 10'h3f2;
        mem[501] = 10'h1d8;
        mem[502] = 10'h31f;
        mem[503] = 10'h35b;
        mem[504] = 10'h100;
        mem[505] = 10'h16b;
        mem[506] = 10'h2e3;
        mem[507] = 10'h1e1;
        mem[508] = 10'h2a4;
        mem[509] = 10'h321;
        mem[510] = 10'h35c;
        mem[511] = 10'h3b3;
        mem[512] = 10'h209;
        mem[513] = 10'h217;
        mem[514] = 10'h361;
        mem[515] = 10'h3d4;
        mem[516] = 10'h120;
        mem[517] = 10'h053;
        mem[518] = 10'h367;
        mem[519] = 10'h20c;
        mem[520] = 10'h398;
        mem[521] = 10'h07e;
        mem[522] = 10'h251;
        mem[523] = 10'h3f6;
        mem[524] = 10'h0cb;
        mem[525] = 10'h25e;
        mem[526] = 10'h2b9;
        mem[527] = 10'h39d;
        mem[528] = 10'h38e;
        mem[529] = 10'h1c6;
        mem[530] = 10'h2dc;
        mem[531] = 10'h1d3;
        mem[532] = 10'h034;
        mem[533] = 10'h272;
        mem[534] = 10'h0db;
        mem[535] = 10'h178;
        mem[536] = 10'h2ed;
        mem[537] = 10'h246;
        mem[538] = 10'h079;
        mem[539] = 10'h098;
        mem[540] = 10'h0b5;
        mem[541] = 10'h0fb;
        mem[542] = 10'h189;
        mem[543] = 10'h078;
        mem[544] = 10'h10c;
        mem[545] = 10'h072;
        mem[546] = 10'h038;
        mem[547] = 10'h1c1;
        mem[548] = 10'h313;
        mem[549] = 10'h3d7;
        mem[550] = 10'h069;
        mem[551] = 10'h1a8;
        mem[552] = 10'h007;
        mem[553] = 10'h16d;
        mem[554] = 10'h2af;
        mem[555] = 10'h317;
        mem[556] = 10'h3f3;
        mem[557] = 10'h101;
        mem[558] = 10'h3ef;
        mem[559] = 10'h262;
        mem[560] = 10'h230;
        mem[561] = 10'h033;
        mem[562] = 10'h1f4;
        mem[563] = 10'h388;
        mem[564] = 10'h04e;
        mem[565] = 10'h311;
        mem[566] = 10'h17e;
        mem[567] = 10'h245;
        mem[568] = 10'h330;
        mem[569] = 10'h0fc;
        mem[570] = 10'h227;
        mem[571] = 10'h2b5;
        mem[572] = 10'h1ac;
        mem[573] = 10'h3ae;
        mem[574] = 10'h3b7;
        mem[575] = 10'h244;
        mem[576] = 10'h3f8;
        mem[577] = 10'h2a3;
        mem[578] = 10'h0a1;
        mem[579] = 10'h350;
        mem[580] = 10'h0b6;
        mem[581] = 10'h1f6;
        mem[582] = 10'h1dc;
        mem[583] = 10'h0da;
        mem[584] = 10'h3bb;
        mem[585] = 10'h0a9;
        mem[586] = 10'h319;
        mem[587] = 10'h10e;
        mem[588] = 10'h3cf;
        mem[589] = 10'h13d;
        mem[590] = 10'h19b;
        mem[591] = 10'h220;
        mem[592] = 10'h29a;
        mem[593] = 10'h12d;
        mem[594] = 10'h0bf;
        mem[595] = 10'h24c;
        mem[596] = 10'h363;
        mem[597] = 10'h0ef;
        mem[598] = 10'h391;
        mem[599] = 10'h0c8;
        mem[600] = 10'h3ce;
        mem[601] = 10'h223;
        mem[602] = 10'h3a8;
        mem[603] = 10'h238;
        mem[604] = 10'h20a;
        mem[605] = 10'h340;
        mem[606] = 10'h15e;
        mem[607] = 10'h060;
        mem[608] = 10'h2d5;
        mem[609] = 10'h284;
        mem[610] = 10'h0ff;
        mem[611] = 10'h2fd;
        mem[612] = 10'h0ab;
        mem[613] = 10'h1e5;
        mem[614] = 10'h1fe;
        mem[615] = 10'h1ab;
        mem[616] = 10'h05f;
        mem[617] = 10'h331;
        mem[618] = 10'h2a2;
        mem[619] = 10'h043;
        mem[620] = 10'h0a8;
        mem[621] = 10'h110;
        mem[622] = 10'h183;
        mem[623] = 10'h028;
        mem[624] = 10'h00d;
        mem[625] = 10'h18b;
        mem[626] = 10'h085;
        mem[627] = 10'h084;
        mem[628] = 10'h25f;
        mem[629] = 10'h0a0;
        mem[630] = 10'h225;
        mem[631] = 10'h3d9;
        mem[632] = 10'h061;
        mem[633] = 10'h045;
        mem[634] = 10'h1cd;
        mem[635] = 10'h1b6;
        mem[636] = 10'h113;
        mem[637] = 10'h28c;
        mem[638] = 10'h3eb;
        mem[639] = 10'h0af;
        mem[640] = 10'h2f1;
        mem[641] = 10'h1f3;
        mem[642] = 10'h0b4;
        mem[643] = 10'h0c2;
        mem[644] = 10'h293;
        mem[645] = 10'h13e;
        mem[646] = 10'h3a9;
        mem[647] = 10'h161;
        mem[648] = 10'h275;
        mem[649] = 10'h1e0;
        mem[650] = 10'h351;
        mem[651] = 10'h0b8;
        mem[652] = 10'h318;
        mem[653] = 10'h150;
        mem[654] = 10'h3e8;
        mem[655] = 10'h2c3;
        mem[656] = 10'h25a;
        mem[657] = 10'h30b;
        mem[658] = 10'h2bb;
        mem[659] = 10'h19c;
        mem[660] = 10'h3b1;
        mem[661] = 10'h19a;
        mem[662] = 10'h202;
        mem[663] = 10'h0ee;
        mem[664] = 10'h373;
        mem[665] = 10'h062;
        mem[666] = 10'h1fa;
        mem[667] = 10'h035;
        mem[668] = 10'h16e;
        mem[669] = 10'h0cf;
        mem[670] = 10'h23d;
        mem[671] = 10'h380;
        mem[672] = 10'h2d1;
        mem[673] = 10'h2cf;
        mem[674] = 10'h17a;
        mem[675] = 10'h2db;
        mem[676] = 10'h397;
        mem[677] = 10'h308;
        mem[678] = 10'h36f;
        mem[679] = 10'h32f;
        mem[680] = 10'h174;
        mem[681] = 10'h38f;
        mem[682] = 10'h3dc;
        mem[683] = 10'h040;
        mem[684] = 10'h121;
        mem[685] = 10'h197;
        mem[686] = 10'h360;
        mem[687] = 10'h05d;
        mem[688] = 10'h04c;
        mem[689] = 10'h126;
        mem[690] = 10'h21d;
        mem[691] = 10'h148;
        mem[692] = 10'h236;
        mem[693] = 10'h3a7;
        mem[694] = 10'h029;
        mem[695] = 10'h010;
        mem[696] = 10'h190;
        mem[697] = 10'h02c;
        mem[698] = 10'h02f;
        mem[699] = 10'h2ec;
        mem[700] = 10'h2d9;
        mem[701] = 10'h29c;
        mem[702] = 10'h31d;
        mem[703] = 10'h222;
        mem[704] = 10'h302;
        mem[705] = 10'h1b2;
        mem[706] = 10'h116;
        mem[707] = 10'h37a;
        mem[708] = 10'h134;
        mem[709] = 10'h3b9;
        mem[710] = 10'h2d2;
        mem[711] = 10'h2b0;
        mem[712] = 10'h0d6;
        mem[713] = 10'h025;
        mem[714] = 10'h1b1;
        mem[715] = 10'h2ea;
        mem[716] = 10'h362;
        mem[717] = 10'h26d;
        mem[718] = 10'h390;
        mem[719] = 10'h24d;
        mem[720] = 10'h35d;
        mem[721] = 10'h173;
        mem[722] = 10'h325;
        mem[723] = 10'h324;
        mem[724] = 10'h28d;
        mem[725] = 10'h2df;
        mem[726] = 10'h285;
        mem[727] = 10'h0c6;
        mem[728] = 10'h39e;
        mem[729] = 10'h2b6;
        mem[730] = 10'h3f7;
        mem[731] = 10'h063;
        mem[732] = 10'h3cd;
        mem[733] = 10'h04d;
        mem[734] = 10'h393;
        mem[735] = 10'h2bf;
        mem[736] = 10'h090;
        mem[737] = 10'h163;
        mem[738] = 10'h0bd;
        mem[739] = 10'h03a;
        mem[740] = 10'h059;
        mem[741] = 10'h19f;
        mem[742] = 10'h1ef;
        mem[743] = 10'h168;
        mem[744] = 10'h287;
        mem[745] = 10'h3c9;
        mem[746] = 10'h1e3;
        mem[747] = 10'h1b0;
        mem[748] = 10'h38c;
        mem[749] = 10'h2a5;
        mem[750] = 10'h1e6;
        mem[751] = 10'h082;
        mem[752] = 10'h051;
        mem[753] = 10'h2f2;
        mem[754] = 10'h344;
        mem[755] = 10'h1ba;
        mem[756] = 10'h3e6;
        mem[757] = 10'h0c1;
        mem[758] = 10'h382;
        mem[759] = 10'h20f;
        mem[760] = 10'h0a5;
        mem[761] = 10'h1bd;
        mem[762] = 10'h097;
        mem[763] = 10'h140;
        mem[764] = 10'h3c6;
        mem[765] = 10'h1cf;
        mem[766] = 10'h369;
        mem[767] = 10'h21a;
        mem[768] = 10'h2e0;
        mem[769] = 10'h096;
        mem[770] = 10'h158;
        mem[771] = 10'h24a;
        mem[772] = 10'h198;
        mem[773] = 10'h179;
        mem[774] = 10'h26f;
        mem[775] = 10'h171;
        mem[776] = 10'h14d;
        mem[777] = 10'h013;
        mem[778] = 10'h306;
        mem[779] = 10'h0c0;
        mem[780] = 10'h349;
        mem[781] = 10'h2e6;
        mem[782] = 10'h207;
        mem[783] = 10'h2b8;
        mem[784] = 10'h12b;
        mem[785] = 10'h254;
        mem[786] = 10'h081;
        mem[787] = 10'h002;
        mem[788] = 10'h288;
        mem[789] = 10'h3a6;
        mem[790] = 10'h001;
        mem[791] = 10'h32b;
        mem[792] = 10'h0f5;
        mem[793] = 10'h337;
        mem[794] = 10'h066;
        mem[795] = 10'h3a5;
        mem[796] = 10'h144;
        mem[797] = 10'h1e9;
        mem[798] = 10'h15b;
        mem[799] = 10'h030;
        mem[800] = 10'h153;
        mem[801] = 10'h102;
        mem[802] = 10'h30c;
        mem[803] = 10'h136;
        mem[804] = 10'h124;
        mem[805] = 10'h019;
        mem[806] = 10'h08c;
        mem[807] = 10'h273;
        mem[808] = 10'h1d2;
        mem[809] = 10'h162;
        mem[810] = 10'h3e1;
        mem[811] = 10'h133;
        mem[812] = 10'h212;
        mem[813] = 10'h290;
        mem[814] = 10'h180;
        mem[815] = 10'h0d9;
        mem[816] = 10'h09c;
        mem[817] = 10'h000;
        mem[818] = 10'h138;
        mem[819] = 10'h14c;
        mem[820] = 10'h135;
        mem[821] = 10'h068;
        mem[822] = 10'h07a;
        mem[823] = 10'h22c;
        mem[824] = 10'h279;
        mem[825] = 10'h268;
        mem[826] = 10'h36a;
        mem[827] = 10'h0bc;
        mem[828] = 10'h3de;
        mem[829] = 10'h228;
        mem[830] = 10'h141;
        mem[831] = 10'h0ec;
        mem[832] = 10'h0aa;
        mem[833] = 10'h235;
        mem[834] = 10'h10f;
        mem[835] = 10'h291;
        mem[836] = 10'h36b;
        mem[837] = 10'h18c;
        mem[838] = 10'h1f1;
        mem[839] = 10'h1be;
        mem[840] = 10'h371;
        mem[841] = 10'h1d0;
        mem[842] = 10'h0e7;
        mem[843] = 10'h37e;
        mem[844] = 10'h248;
        mem[845] = 10'h24b;
        mem[846] = 10'h26e;
        mem[847] = 10'h395;
        mem[848] = 10'h1ec;
        mem[849] = 10'h21b;
        mem[850] = 10'h358;
        mem[851] = 10'h277;
        mem[852] = 10'h19e;
        mem[853] = 10'h2c8;
        mem[854] = 10'h19d;
        mem[855] = 10'h194;
        mem[856] = 10'h341;
        mem[857] = 10'h259;
        mem[858] = 10'h2f8;
        mem[859] = 10'h023;
        mem[860] = 10'h039;
        mem[861] = 10'h151;
        mem[862] = 10'h39c;
        mem[863] = 10'h3bc;
        mem[864] = 10'h3fe;
        mem[865] = 10'h0a4;
        mem[866] = 10'h2cc;
        mem[867] = 10'h1ea;
        mem[868] = 10'h06a;
        mem[869] = 10'h02d;
        mem[870] = 10'h0b1;
        mem[871] = 10'h08d;
        mem[872] = 10'h1d4;
        mem[873] = 10'h055;
        mem[874] = 10'h03e;
        mem[875] = 10'h00b;
        mem[876] = 10'h267;
        mem[877] = 10'h01d;
        mem[878] = 10'h0df;
        mem[879] = 10'h160;
        mem[880] = 10'h10a;
        mem[881] = 10'h157;
        mem[882] = 10'h1b3;
        mem[883] = 10'h21e;
        mem[884] = 10'h155;
        mem[885] = 10'h0ac;
        mem[886] = 10'h30f;
        mem[887] = 10'h1b9;
        mem[888] = 10'h0b2;
        mem[889] = 10'h224;
        mem[890] = 10'h334;
        mem[891] = 10'h214;
        mem[892] = 10'h065;
        mem[893] = 10'h165;
        mem[894] = 10'h366;
        mem[895] = 10'h323;
        mem[896] = 10'h274;
        mem[897] = 10'h39f;
        mem[898] = 10'h3af;
        mem[899] = 10'h12c;
        mem[900] = 10'h094;
        mem[901] = 10'h074;
        mem[902] = 10'h105;
        mem[903] = 10'h0ca;
        mem[904] = 10'h1d6;
        mem[905] = 10'h381;
        mem[906] = 10'h087;
        mem[907] = 10'h15a;
        mem[908] = 10'h17c;
        mem[909] = 10'h3c0;
        mem[910] = 10'h004;
        mem[911] = 10'h29f;
        mem[912] = 10'h234;
        mem[913] = 10'h2f5;
        mem[914] = 10'h14a;
        mem[915] = 10'h3b6;
        mem[916] = 10'h25b;
        mem[917] = 10'h2eb;
        mem[918] = 10'h22b;
        mem[919] = 10'h12e;
        mem[920] = 10'h2de;
        mem[921] = 10'h34b;
        mem[922] = 10'h24e;
        mem[923] = 10'h2e7;
        mem[924] = 10'h3c3;
        mem[925] = 10'h233;
        mem[926] = 10'h003;
        mem[927] = 10'h345;
        mem[928] = 10'h260;
        mem[929] = 10'h064;
        mem[930] = 10'h23a;
        mem[931] = 10'h356;
        mem[932] = 10'h18d;
        mem[933] = 10'h2fb;
        mem[934] = 10'h22d;
        mem[935] = 10'h34a;
        mem[936] = 10'h27b;
        mem[937] = 10'h130;
        mem[938] = 10'h243;
        mem[939] = 10'h077;
        mem[940] = 10'h38a;
        mem[941] = 10'h12a;
        mem[942] = 10'h091;
        mem[943] = 10'h103;
        mem[944] = 10'h21f;
        mem[945] = 10'h1f2;
        mem[946] = 10'h09d;
        mem[947] = 10'h009;
        mem[948] = 10'h16f;
        mem[949] = 10'h396;
        mem[950] = 10'h3a3;
        mem[951] = 10'h0be;
        mem[952] = 10'h376;
        mem[953] = 10'h2f6;
        mem[954] = 10'h2a7;
        mem[955] = 10'h067;
        mem[956] = 10'h339;
        mem[957] = 10'h27d;
        mem[958] = 10'h377;
        mem[959] = 10'h2e2;
        mem[960] = 10'h1e2;
        mem[961] = 10'h263;
        mem[962] = 10'h29e;
        mem[963] = 10'h39a;
        mem[964] = 10'h1bb;
        mem[965] = 10'h3b5;
        mem[966] = 10'h156;
        mem[967] = 10'h22f;
        mem[968] = 10'h3ca;
        mem[969] = 10'h3ed;
        mem[970] = 10'h128;
        mem[971] = 10'h070;
        mem[972] = 10'h1e8;
        mem[973] = 10'h1a5;
        mem[974] = 10'h3fa;
        mem[975] = 10'h09a;
        mem[976] = 10'h252;
        mem[977] = 10'h118;
        mem[978] = 10'h33d;
        mem[979] = 10'h20e;
        mem[980] = 10'h1df;
        mem[981] = 10'h131;
        mem[982] = 10'h309;
        mem[983] = 10'h107;
        mem[984] = 10'h33b;
        mem[985] = 10'h047;
        mem[986] = 10'h229;
        mem[987] = 10'h37f;
        mem[988] = 10'h1ed;
        mem[989] = 10'h30a;
        mem[990] = 10'h3d5;
        mem[991] = 10'h0b9;
        mem[992] = 10'h09f;
        mem[993] = 10'h02b;
        mem[994] = 10'h3f9;
        mem[995] = 10'h28b;
        mem[996] = 10'h05a;
        mem[997] = 10'h241;
        mem[998] = 10'h1fb;
        mem[999] = 10'h266;
        mem[1000] = 10'h184;
        mem[1001] = 10'h108;
        mem[1002] = 10'h16c;
        mem[1003] = 10'h384;
        mem[1004] = 10'h270;
        mem[1005] = 10'h170;
        mem[1006] = 10'h399;
        mem[1007] = 10'h3c7;
        mem[1008] = 10'h10d;
        mem[1009] = 10'h11e;
        mem[1010] = 10'h193;
        mem[1011] = 10'h0b7;
        mem[1012] = 10'h322;
        mem[1013] = 10'h298;
        mem[1014] = 10'h075;
        mem[1015] = 10'h336;
        mem[1016] = 10'h02a;
        mem[1017] = 10'h208;
        mem[1018] = 10'h042;
        mem[1019] = 10'h2ef;
        mem[1020] = 10'h27c;
        mem[1021] = 10'h2d6;
        mem[1022] = 10'h3a4;
        mem[1023] = 10'h3f4;
    end
endmodule

module encrypt_4sbox_large2(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h0a1;
        mem[1] = 10'h315;
        mem[2] = 10'h066;
        mem[3] = 10'h0a4;
        mem[4] = 10'h0bc;
        mem[5] = 10'h0bd;
        mem[6] = 10'h3b0;
        mem[7] = 10'h248;
        mem[8] = 10'h095;
        mem[9] = 10'h24f;
        mem[10] = 10'h073;
        mem[11] = 10'h025;
        mem[12] = 10'h0f0;
        mem[13] = 10'h053;
        mem[14] = 10'h1ec;
        mem[15] = 10'h3ac;
        mem[16] = 10'h394;
        mem[17] = 10'h2d8;
        mem[18] = 10'h187;
        mem[19] = 10'h02d;
        mem[20] = 10'h299;
        mem[21] = 10'h3ad;
        mem[22] = 10'h273;
        mem[23] = 10'h3c1;
        mem[24] = 10'h139;
        mem[25] = 10'h077;
        mem[26] = 10'h2f1;
        mem[27] = 10'h07d;
        mem[28] = 10'h284;
        mem[29] = 10'h03b;
        mem[30] = 10'h1d4;
        mem[31] = 10'h3e7;
        mem[32] = 10'h316;
        mem[33] = 10'h136;
        mem[34] = 10'h293;
        mem[35] = 10'h3cc;
        mem[36] = 10'h1ce;
        mem[37] = 10'h19f;
        mem[38] = 10'h17c;
        mem[39] = 10'h048;
        mem[40] = 10'h201;
        mem[41] = 10'h18b;
        mem[42] = 10'h22b;
        mem[43] = 10'h0a2;
        mem[44] = 10'h2c2;
        mem[45] = 10'h267;
        mem[46] = 10'h265;
        mem[47] = 10'h308;
        mem[48] = 10'h0fe;
        mem[49] = 10'h208;
        mem[50] = 10'h3e6;
        mem[51] = 10'h2f4;
        mem[52] = 10'h256;
        mem[53] = 10'h110;
        mem[54] = 10'h13b;
        mem[55] = 10'h156;
        mem[56] = 10'h1b8;
        mem[57] = 10'h11b;
        mem[58] = 10'h32b;
        mem[59] = 10'h2ee;
        mem[60] = 10'h3d8;
        mem[61] = 10'h22e;
        mem[62] = 10'h125;
        mem[63] = 10'h1ee;
        mem[64] = 10'h28f;
        mem[65] = 10'h2a9;
        mem[66] = 10'h38c;
        mem[67] = 10'h33f;
        mem[68] = 10'h289;
        mem[69] = 10'h266;
        mem[70] = 10'h1fd;
        mem[71] = 10'h21b;
        mem[72] = 10'h1fe;
        mem[73] = 10'h26d;
        mem[74] = 10'h2a3;
        mem[75] = 10'h3ed;
        mem[76] = 10'h36e;
        mem[77] = 10'h2f7;
        mem[78] = 10'h32f;
        mem[79] = 10'h3c6;
        mem[80] = 10'h211;
        mem[81] = 10'h301;
        mem[82] = 10'h383;
        mem[83] = 10'h10d;
        mem[84] = 10'h1a1;
        mem[85] = 10'h166;
        mem[86] = 10'h0bf;
        mem[87] = 10'h2b2;
        mem[88] = 10'h10a;
        mem[89] = 10'h028;
        mem[90] = 10'h291;
        mem[91] = 10'h216;
        mem[92] = 10'h241;
        mem[93] = 10'h097;
        mem[94] = 10'h05c;
        mem[95] = 10'h3ee;
        mem[96] = 10'h006;
        mem[97] = 10'h1e9;
        mem[98] = 10'h3fc;
        mem[99] = 10'h19e;
        mem[100] = 10'h051;
        mem[101] = 10'h1e5;
        mem[102] = 10'h0ed;
        mem[103] = 10'h381;
        mem[104] = 10'h043;
        mem[105] = 10'h0e1;
        mem[106] = 10'h275;
        mem[107] = 10'h005;
        mem[108] = 10'h23a;
        mem[109] = 10'h2bc;
        mem[110] = 10'h29b;
        mem[111] = 10'h2d0;
        mem[112] = 10'h3a0;
        mem[113] = 10'h240;
        mem[114] = 10'h0a5;
        mem[115] = 10'h2b1;
        mem[116] = 10'h217;
        mem[117] = 10'h0e3;
        mem[118] = 10'h05f;
        mem[119] = 10'h15d;
        mem[120] = 10'h35c;
        mem[121] = 10'h12e;
        mem[122] = 10'h1b1;
        mem[123] = 10'h3f3;
        mem[124] = 10'h2fe;
        mem[125] = 10'h30d;
        mem[126] = 10'h1a5;
        mem[127] = 10'h108;
        mem[128] = 10'h399;
        mem[129] = 10'h332;
        mem[130] = 10'h27e;
        mem[131] = 10'h03e;
        mem[132] = 10'h304;
        mem[133] = 10'h2c9;
        mem[134] = 10'h20f;
        mem[135] = 10'h163;
        mem[136] = 10'h0f3;
        mem[137] = 10'h3a1;
        mem[138] = 10'h378;
        mem[139] = 10'h395;
        mem[140] = 10'h1ff;
        mem[141] = 10'h0d9;
        mem[142] = 10'h24e;
        mem[143] = 10'h2e9;
        mem[144] = 10'h2c4;
        mem[145] = 10'h328;
        mem[146] = 10'h0fb;
        mem[147] = 10'h339;
        mem[148] = 10'h0b8;
        mem[149] = 10'h281;
        mem[150] = 10'h14a;
        mem[151] = 10'h03a;
        mem[152] = 10'h2bd;
        mem[153] = 10'h325;
        mem[154] = 10'h385;
        mem[155] = 10'h175;
        mem[156] = 10'h21f;
        mem[157] = 10'h17e;
        mem[158] = 10'h232;
        mem[159] = 10'h3d4;
        mem[160] = 10'h052;
        mem[161] = 10'h26a;
        mem[162] = 10'h29a;
        mem[163] = 10'h19a;
        mem[164] = 10'h2bf;
        mem[165] = 10'h340;
        mem[166] = 10'h15b;
        mem[167] = 10'h38f;
        mem[168] = 10'h311;
        mem[169] = 10'h288;
        mem[170] = 10'h398;
        mem[171] = 10'h2e0;
        mem[172] = 10'h396;
        mem[173] = 10'h20e;
        mem[174] = 10'h138;
        mem[175] = 10'h1be;
        mem[176] = 10'h0ab;
        mem[177] = 10'h19d;
        mem[178] = 10'h3ea;
        mem[179] = 10'h1ac;
        mem[180] = 10'h359;
        mem[181] = 10'h007;
        mem[182] = 10'h0c6;
        mem[183] = 10'h302;
        mem[184] = 10'h2a1;
        mem[185] = 10'h274;
        mem[186] = 10'h3e5;
        mem[187] = 10'h12a;
        mem[188] = 10'h24d;
        mem[189] = 10'h295;
        mem[190] = 10'h0c4;
        mem[191] = 10'h04d;
        mem[192] = 10'h37c;
        mem[193] = 10'h3c2;
        mem[194] = 10'h21d;
        mem[195] = 10'h3db;
        mem[196] = 10'h2ea;
        mem[197] = 10'h1ab;
        mem[198] = 10'h05b;
        mem[199] = 10'h01a;
        mem[200] = 10'h150;
        mem[201] = 10'h1d3;
        mem[202] = 10'h2f3;
        mem[203] = 10'h0ef;
        mem[204] = 10'h182;
        mem[205] = 10'h1bf;
        mem[206] = 10'h16d;
        mem[207] = 10'h29f;
        mem[208] = 10'h37f;
        mem[209] = 10'h39b;
        mem[210] = 10'h2ef;
        mem[211] = 10'h36a;
        mem[212] = 10'h019;
        mem[213] = 10'h3a5;
        mem[214] = 10'h1f2;
        mem[215] = 10'h1f1;
        mem[216] = 10'h104;
        mem[217] = 10'h12b;
        mem[218] = 10'h1bc;
        mem[219] = 10'h34e;
        mem[220] = 10'h01b;
        mem[221] = 10'h002;
        mem[222] = 10'h1a3;
        mem[223] = 10'h0a9;
        mem[224] = 10'h098;
        mem[225] = 10'h031;
        mem[226] = 10'h1f8;
        mem[227] = 10'h1af;
        mem[228] = 10'h3a3;
        mem[229] = 10'h176;
        mem[230] = 10'h247;
        mem[231] = 10'h249;
        mem[232] = 10'h33b;
        mem[233] = 10'h13d;
        mem[234] = 10'h314;
        mem[235] = 10'h366;
        mem[236] = 10'h35f;
        mem[237] = 10'h254;
        mem[238] = 10'h319;
        mem[239] = 10'h3af;
        mem[240] = 10'h0cd;
        mem[241] = 10'h02a;
        mem[242] = 10'h2b7;
        mem[243] = 10'h04b;
        mem[244] = 10'h0a3;
        mem[245] = 10'h068;
        mem[246] = 10'h1b0;
        mem[247] = 10'h03f;
        mem[248] = 10'h320;
        mem[249] = 10'h19b;
        mem[250] = 10'h337;
        mem[251] = 10'h2cb;
        mem[252] = 10'h3d6;
        mem[253] = 10'h2e8;
        mem[254] = 10'h338;
        mem[255] = 10'h259;
        mem[256] = 10'h2cf;
        mem[257] = 10'h32a;
        mem[258] = 10'h107;
        mem[259] = 10'h00c;
        mem[260] = 10'h1c4;
        mem[261] = 10'h10b;
        mem[262] = 10'h16b;
        mem[263] = 10'h056;
        mem[264] = 10'h1b5;
        mem[265] = 10'h10e;
        mem[266] = 10'h27c;
        mem[267] = 10'h0bb;
        mem[268] = 10'h357;
        mem[269] = 10'h34f;
        mem[270] = 10'h3b5;
        mem[271] = 10'h25a;
        mem[272] = 10'h197;
        mem[273] = 10'h0ee;
        mem[274] = 10'h022;
        mem[275] = 10'h015;
        mem[276] = 10'h1c9;
        mem[277] = 10'h1e1;
        mem[278] = 10'h08c;
        mem[279] = 10'h3da;
        mem[280] = 10'h341;
        mem[281] = 10'h059;
        mem[282] = 10'h348;
        mem[283] = 10'h3b9;
        mem[284] = 10'h218;
        mem[285] = 10'h2ce;
        mem[286] = 10'h1f5;
        mem[287] = 10'h21c;
        mem[288] = 10'h2d1;
        mem[289] = 10'h23f;
        mem[290] = 10'h3ce;
        mem[291] = 10'h061;
        mem[292] = 10'h3a4;
        mem[293] = 10'h135;
        mem[294] = 10'h3c8;
        mem[295] = 10'h212;
        mem[296] = 10'h16c;
        mem[297] = 10'h2df;
        mem[298] = 10'h283;
        mem[299] = 10'h28b;
        mem[300] = 10'h252;
        mem[301] = 10'h121;
        mem[302] = 10'h23c;
        mem[303] = 10'h38a;
        mem[304] = 10'h2b8;
        mem[305] = 10'h228;
        mem[306] = 10'h055;
        mem[307] = 10'h2a6;
        mem[308] = 10'h195;
        mem[309] = 10'h3aa;
        mem[310] = 10'h2a5;
        mem[311] = 10'h06b;
        mem[312] = 10'h3a7;
        mem[313] = 10'h37b;
        mem[314] = 10'h243;
        mem[315] = 10'h39d;
        mem[316] = 10'h038;
        mem[317] = 10'h257;
        mem[318] = 10'h36f;
        mem[319] = 10'h321;
        mem[320] = 10'h3c5;
        mem[321] = 10'h0d6;
        mem[322] = 10'h371;
        mem[323] = 10'h268;
        mem[324] = 10'h1ed;
        mem[325] = 10'h1f3;
        mem[326] = 10'h36b;
        mem[327] = 10'h191;
        mem[328] = 10'h167;
        mem[329] = 10'h296;
        mem[330] = 10'h0d0;
        mem[331] = 10'h189;
        mem[332] = 10'h1a4;
        mem[333] = 10'h089;
        mem[334] = 10'h392;
        mem[335] = 10'h3d7;
        mem[336] = 10'h2ff;
        mem[337] = 10'h072;
        mem[338] = 10'h346;
        mem[339] = 10'h30b;
        mem[340] = 10'h04a;
        mem[341] = 10'h188;
        mem[342] = 10'h16a;
        mem[343] = 10'h1d5;
        mem[344] = 10'h313;
        mem[345] = 10'h202;
        mem[346] = 10'h356;
        mem[347] = 10'h2d4;
        mem[348] = 10'h3c9;
        mem[349] = 10'h306;
        mem[350] = 10'h016;
        mem[351] = 10'h2ac;
        mem[352] = 10'h37e;
        mem[353] = 10'h3b2;
        mem[354] = 10'h207;
        mem[355] = 10'h2a4;
        mem[356] = 10'h269;
        mem[357] = 10'h02e;
        mem[358] = 10'h361;
        mem[359] = 10'h226;
        mem[360] = 10'h303;
        mem[361] = 10'h181;
        mem[362] = 10'h079;
        mem[363] = 10'h1c3;
        mem[364] = 10'h1b9;
        mem[365] = 10'h0dc;
        mem[366] = 10'h001;
        mem[367] = 10'h129;
        mem[368] = 10'h33a;
        mem[369] = 10'h1b3;
        mem[370] = 10'h01e;
        mem[371] = 10'h344;
        mem[372] = 10'h09a;
        mem[373] = 10'h0d3;
        mem[374] = 10'h2c0;
        mem[375] = 10'h264;
        mem[376] = 10'h100;
        mem[377] = 10'h3f6;
        mem[378] = 10'h17d;
        mem[379] = 10'h041;
        mem[380] = 10'h1b4;
        mem[381] = 10'h0af;
        mem[382] = 10'h3b8;
        mem[383] = 10'h387;
        mem[384] = 10'h2d3;
        mem[385] = 10'h3e8;
        mem[386] = 10'h0eb;
        mem[387] = 10'h376;
        mem[388] = 10'h1f9;
        mem[389] = 10'h071;
        mem[390] = 10'h285;
        mem[391] = 10'h27b;
        mem[392] = 10'h07e;
        mem[393] = 10'h145;
        mem[394] = 10'h02c;
        mem[395] = 10'h09b;
        mem[396] = 10'h040;
        mem[397] = 10'h238;
        mem[398] = 10'h389;
        mem[399] = 10'h021;
        mem[400] = 10'h298;
        mem[401] = 10'h20a;
        mem[402] = 10'h20d;
        mem[403] = 10'h300;
        mem[404] = 10'h113;
        mem[405] = 10'h377;
        mem[406] = 10'h31d;
        mem[407] = 10'h26c;
        mem[408] = 10'h33c;
        mem[409] = 10'h0c5;
        mem[410] = 10'h3df;
        mem[411] = 10'h0d2;
        mem[412] = 10'h1d9;
        mem[413] = 10'h04c;
        mem[414] = 10'h276;
        mem[415] = 10'h1fb;
        mem[416] = 10'h0b4;
        mem[417] = 10'h2cc;
        mem[418] = 10'h023;
        mem[419] = 10'h08e;
        mem[420] = 10'h2d9;
        mem[421] = 10'h27d;
        mem[422] = 10'h364;
        mem[423] = 10'h3fe;
        mem[424] = 10'h199;
        mem[425] = 10'h2ae;
        mem[426] = 10'h32d;
        mem[427] = 10'h15c;
        mem[428] = 10'h0a7;
        mem[429] = 10'h034;
        mem[430] = 10'h06d;
        mem[431] = 10'h117;
        mem[432] = 10'h06c;
        mem[433] = 10'h03c;
        mem[434] = 10'h3d5;
        mem[435] = 10'h37d;
        mem[436] = 10'h101;
        mem[437] = 10'h1ba;
        mem[438] = 10'h103;
        mem[439] = 10'h137;
        mem[440] = 10'h198;
        mem[441] = 10'h28e;
        mem[442] = 10'h00f;
        mem[443] = 10'h143;
        mem[444] = 10'h08d;
        mem[445] = 10'h1f0;
        mem[446] = 10'h33e;
        mem[447] = 10'h35b;
        mem[448] = 10'h000;
        mem[449] = 10'h30f;
        mem[450] = 10'h260;
        mem[451] = 10'h004;
        mem[452] = 10'h20b;
        mem[453] = 10'h0f5;
        mem[454] = 10'h0f1;
        mem[455] = 10'h3d3;
        mem[456] = 10'h0b3;
        mem[457] = 10'h0f7;
        mem[458] = 10'h084;
        mem[459] = 10'h2f6;
        mem[460] = 10'h32c;
        mem[461] = 10'h258;
        mem[462] = 10'h036;
        mem[463] = 10'h0ad;
        mem[464] = 10'h2be;
        mem[465] = 10'h109;
        mem[466] = 10'h230;
        mem[467] = 10'h00e;
        mem[468] = 10'h305;
        mem[469] = 10'h2e3;
        mem[470] = 10'h09d;
        mem[471] = 10'h179;
        mem[472] = 10'h270;
        mem[473] = 10'h229;
        mem[474] = 10'h050;
        mem[475] = 10'h224;
        mem[476] = 10'h2e6;
        mem[477] = 10'h127;
        mem[478] = 10'h2cd;
        mem[479] = 10'h1fa;
        mem[480] = 10'h1a0;
        mem[481] = 10'h1de;
        mem[482] = 10'h3fa;
        mem[483] = 10'h058;
        mem[484] = 10'h0da;
        mem[485] = 10'h204;
        mem[486] = 10'h119;
        mem[487] = 10'h123;
        mem[488] = 10'h2eb;
        mem[489] = 10'h33d;
        mem[490] = 10'h326;
        mem[491] = 10'h203;
        mem[492] = 10'h244;
        mem[493] = 10'h07f;
        mem[494] = 10'h39a;
        mem[495] = 10'h331;
        mem[496] = 10'h362;
        mem[497] = 10'h0d1;
        mem[498] = 10'h0c8;
        mem[499] = 10'h148;
        mem[500] = 10'h1c8;
        mem[501] = 10'h3ba;
        mem[502] = 10'h014;
        mem[503] = 10'h069;
        mem[504] = 10'h292;
        mem[505] = 10'h375;
        mem[506] = 10'h3d0;
        mem[507] = 10'h358;
        mem[508] = 10'h196;
        mem[509] = 10'h286;
        mem[510] = 10'h12f;
        mem[511] = 10'h3dc;
        mem[512] = 10'h102;
        mem[513] = 10'h14f;
        mem[514] = 10'h1c6;
        mem[515] = 10'h012;
        mem[516] = 10'h365;
        mem[517] = 10'h1a8;
        mem[518] = 10'h132;
        mem[519] = 10'h38e;
        mem[520] = 10'h01d;
        mem[521] = 10'h367;
        mem[522] = 10'h2aa;
        mem[523] = 10'h39e;
        mem[524] = 10'h2bb;
        mem[525] = 10'h310;
        mem[526] = 10'h1f6;
        mem[527] = 10'h134;
        mem[528] = 10'h146;
        mem[529] = 10'h044;
        mem[530] = 10'h0c3;
        mem[531] = 10'h153;
        mem[532] = 10'h0f4;
        mem[533] = 10'h390;
        mem[534] = 10'h0e7;
        mem[535] = 10'h379;
        mem[536] = 10'h064;
        mem[537] = 10'h215;
        mem[538] = 10'h24a;
        mem[539] = 10'h1a9;
        mem[540] = 10'h12c;
        mem[541] = 10'h206;
        mem[542] = 10'h277;
        mem[543] = 10'h116;
        mem[544] = 10'h3eb;
        mem[545] = 10'h2a8;
        mem[546] = 10'h2fd;
        mem[547] = 10'h08f;
        mem[548] = 10'h06a;
        mem[549] = 10'h05a;
        mem[550] = 10'h2f0;
        mem[551] = 10'h1e8;
        mem[552] = 10'h1d2;
        mem[553] = 10'h30e;
        mem[554] = 10'h29c;
        mem[555] = 10'h0e0;
        mem[556] = 10'h1a7;
        mem[557] = 10'h0fc;
        mem[558] = 10'h3de;
        mem[559] = 10'h1b7;
        mem[560] = 10'h22d;
        mem[561] = 10'h154;
        mem[562] = 10'h30c;
        mem[563] = 10'h3e3;
        mem[564] = 10'h2f9;
        mem[565] = 10'h027;
        mem[566] = 10'h2b4;
        mem[567] = 10'h278;
        mem[568] = 10'h38b;
        mem[569] = 10'h330;
        mem[570] = 10'h0a0;
        mem[571] = 10'h13f;
        mem[572] = 10'h01f;
        mem[573] = 10'h246;
        mem[574] = 10'h0e2;
        mem[575] = 10'h054;
        mem[576] = 10'h29d;
        mem[577] = 10'h2e5;
        mem[578] = 10'h262;
        mem[579] = 10'h21e;
        mem[580] = 10'h347;
        mem[581] = 10'h1b6;
        mem[582] = 10'h169;
        mem[583] = 10'h0ea;
        mem[584] = 10'h082;
        mem[585] = 10'h2c5;
        mem[586] = 10'h180;
        mem[587] = 10'h1b2;
        mem[588] = 10'h070;
        mem[589] = 10'h3bb;
        mem[590] = 10'h350;
        mem[591] = 10'h2ec;
        mem[592] = 10'h030;
        mem[593] = 10'h18c;
        mem[594] = 10'h1fc;
        mem[595] = 10'h2f2;
        mem[596] = 10'h083;
        mem[597] = 10'h11c;
        mem[598] = 10'h1ca;
        mem[599] = 10'h297;
        mem[600] = 10'h0be;
        mem[601] = 10'h28a;
        mem[602] = 10'h200;
        mem[603] = 10'h00d;
        mem[604] = 10'h093;
        mem[605] = 10'h0dd;
        mem[606] = 10'h09c;
        mem[607] = 10'h2a2;
        mem[608] = 10'h236;
        mem[609] = 10'h3ec;
        mem[610] = 10'h0d4;
        mem[611] = 10'h2d2;
        mem[612] = 10'h164;
        mem[613] = 10'h11f;
        mem[614] = 10'h317;
        mem[615] = 10'h2b0;
        mem[616] = 10'h3f0;
        mem[617] = 10'h178;
        mem[618] = 10'h126;
        mem[619] = 10'h057;
        mem[620] = 10'h16e;
        mem[621] = 10'h09e;
        mem[622] = 10'h0e5;
        mem[623] = 10'h1dd;
        mem[624] = 10'h272;
        mem[625] = 10'h234;
        mem[626] = 10'h3d9;
        mem[627] = 10'h34d;
        mem[628] = 10'h149;
        mem[629] = 10'h07c;
        mem[630] = 10'h345;
        mem[631] = 10'h075;
        mem[632] = 10'h3b7;
        mem[633] = 10'h2b6;
        mem[634] = 10'h122;
        mem[635] = 10'h353;
        mem[636] = 10'h076;
        mem[637] = 10'h322;
        mem[638] = 10'h2e4;
        mem[639] = 10'h2c1;
        mem[640] = 10'h1ae;
        mem[641] = 10'h2e2;
        mem[642] = 10'h27a;
        mem[643] = 10'h133;
        mem[644] = 10'h29e;
        mem[645] = 10'h14b;
        mem[646] = 10'h329;
        mem[647] = 10'h1cf;
        mem[648] = 10'h2b5;
        mem[649] = 10'h010;
        mem[650] = 10'h391;
        mem[651] = 10'h25c;
        mem[652] = 10'h223;
        mem[653] = 10'h374;
        mem[654] = 10'h26e;
        mem[655] = 10'h171;
        mem[656] = 10'h3cd;
        mem[657] = 10'h13c;
        mem[658] = 10'h09f;
        mem[659] = 10'h060;
        mem[660] = 10'h1e6;
        mem[661] = 10'h035;
        mem[662] = 10'h1dc;
        mem[663] = 10'h1c0;
        mem[664] = 10'h354;
        mem[665] = 10'h227;
        mem[666] = 10'h2fa;
        mem[667] = 10'h0b6;
        mem[668] = 10'h094;
        mem[669] = 10'h151;
        mem[670] = 10'h324;
        mem[671] = 10'h209;
        mem[672] = 10'h074;
        mem[673] = 10'h3cf;
        mem[674] = 10'h065;
        mem[675] = 10'h213;
        mem[676] = 10'h0cf;
        mem[677] = 10'h307;
        mem[678] = 10'h1cc;
        mem[679] = 10'h063;
        mem[680] = 10'h0b5;
        mem[681] = 10'h1bd;
        mem[682] = 10'h162;
        mem[683] = 10'h237;
        mem[684] = 10'h3be;
        mem[685] = 10'h032;
        mem[686] = 10'h2db;
        mem[687] = 10'h13a;
        mem[688] = 10'h214;
        mem[689] = 10'h0ae;
        mem[690] = 10'h25d;
        mem[691] = 10'h2d7;
        mem[692] = 10'h155;
        mem[693] = 10'h1e3;
        mem[694] = 10'h28d;
        mem[695] = 10'h020;
        mem[696] = 10'h26b;
        mem[697] = 10'h271;
        mem[698] = 10'h3f8;
        mem[699] = 10'h1a2;
        mem[700] = 10'h0f6;
        mem[701] = 10'h3ae;
        mem[702] = 10'h080;
        mem[703] = 10'h349;
        mem[704] = 10'h173;
        mem[705] = 10'h0a6;
        mem[706] = 10'h12d;
        mem[707] = 10'h3e2;
        mem[708] = 10'h30a;
        mem[709] = 10'h31b;
        mem[710] = 10'h1c7;
        mem[711] = 10'h352;
        mem[712] = 10'h05d;
        mem[713] = 10'h177;
        mem[714] = 10'h34c;
        mem[715] = 10'h290;
        mem[716] = 10'h1d7;
        mem[717] = 10'h1d0;
        mem[718] = 10'h0cb;
        mem[719] = 10'h0ce;
        mem[720] = 10'h205;
        mem[721] = 10'h360;
        mem[722] = 10'h18a;
        mem[723] = 10'h078;
        mem[724] = 10'h013;
        mem[725] = 10'h0a8;
        mem[726] = 10'h21a;
        mem[727] = 10'h2d6;
        mem[728] = 10'h1ea;
        mem[729] = 10'h017;
        mem[730] = 10'h3ff;
        mem[731] = 10'h22a;
        mem[732] = 10'h144;
        mem[733] = 10'h1e4;
        mem[734] = 10'h2ed;
        mem[735] = 10'h253;
        mem[736] = 10'h222;
        mem[737] = 10'h3e0;
        mem[738] = 10'h251;
        mem[739] = 10'h323;
        mem[740] = 10'h06e;
        mem[741] = 10'h1c2;
        mem[742] = 10'h221;
        mem[743] = 10'h3a6;
        mem[744] = 10'h0b9;
        mem[745] = 10'h225;
        mem[746] = 10'h2fb;
        mem[747] = 10'h294;
        mem[748] = 10'h1df;
        mem[749] = 10'h003;
        mem[750] = 10'h147;
        mem[751] = 10'h118;
        mem[752] = 10'h067;
        mem[753] = 10'h2e1;
        mem[754] = 10'h0ec;
        mem[755] = 10'h351;
        mem[756] = 10'h31c;
        mem[757] = 10'h04f;
        mem[758] = 10'h2b9;
        mem[759] = 10'h00b;
        mem[760] = 10'h342;
        mem[761] = 10'h3fd;
        mem[762] = 10'h2c6;
        mem[763] = 10'h086;
        mem[764] = 10'h0ff;
        mem[765] = 10'h05e;
        mem[766] = 10'h369;
        mem[767] = 10'h250;
        mem[768] = 10'h185;
        mem[769] = 10'h029;
        mem[770] = 10'h24b;
        mem[771] = 10'h0c2;
        mem[772] = 10'h393;
        mem[773] = 10'h0b2;
        mem[774] = 10'h105;
        mem[775] = 10'h2dc;
        mem[776] = 10'h2a0;
        mem[777] = 10'h3b6;
        mem[778] = 10'h0d8;
        mem[779] = 10'h1db;
        mem[780] = 10'h2af;
        mem[781] = 10'h0aa;
        mem[782] = 10'h210;
        mem[783] = 10'h39c;
        mem[784] = 10'h34a;
        mem[785] = 10'h158;
        mem[786] = 10'h318;
        mem[787] = 10'h343;
        mem[788] = 10'h161;
        mem[789] = 10'h08b;
        mem[790] = 10'h140;
        mem[791] = 10'h368;
        mem[792] = 10'h0cc;
        mem[793] = 10'h092;
        mem[794] = 10'h327;
        mem[795] = 10'h3f1;
        mem[796] = 10'h168;
        mem[797] = 10'h386;
        mem[798] = 10'h018;
        mem[799] = 10'h1cb;
        mem[800] = 10'h193;
        mem[801] = 10'h114;
        mem[802] = 10'h3fb;
        mem[803] = 10'h14c;
        mem[804] = 10'h3e9;
        mem[805] = 10'h2f5;
        mem[806] = 10'h18d;
        mem[807] = 10'h3f5;
        mem[808] = 10'h026;
        mem[809] = 10'h2c7;
        mem[810] = 10'h1c5;
        mem[811] = 10'h174;
        mem[812] = 10'h141;
        mem[813] = 10'h16f;
        mem[814] = 10'h38d;
        mem[815] = 10'h2b3;
        mem[816] = 10'h152;
        mem[817] = 10'h0e8;
        mem[818] = 10'h0f8;
        mem[819] = 10'h2e7;
        mem[820] = 10'h3f4;
        mem[821] = 10'h0f2;
        mem[822] = 10'h335;
        mem[823] = 10'h2a7;
        mem[824] = 10'h35e;
        mem[825] = 10'h10f;
        mem[826] = 10'h27f;
        mem[827] = 10'h2c8;
        mem[828] = 10'h0e4;
        mem[829] = 10'h087;
        mem[830] = 10'h3c7;
        mem[831] = 10'h1e2;
        mem[832] = 10'h3bd;
        mem[833] = 10'h062;
        mem[834] = 10'h0c7;
        mem[835] = 10'h192;
        mem[836] = 10'h0b0;
        mem[837] = 10'h279;
        mem[838] = 10'h04e;
        mem[839] = 10'h3a2;
        mem[840] = 10'h008;
        mem[841] = 10'h15e;
        mem[842] = 10'h165;
        mem[843] = 10'h309;
        mem[844] = 10'h25e;
        mem[845] = 10'h183;
        mem[846] = 10'h280;
        mem[847] = 10'h0e9;
        mem[848] = 10'h19c;
        mem[849] = 10'h011;
        mem[850] = 10'h085;
        mem[851] = 10'h333;
        mem[852] = 10'h024;
        mem[853] = 10'h088;
        mem[854] = 10'h3d2;
        mem[855] = 10'h20c;
        mem[856] = 10'h334;
        mem[857] = 10'h26f;
        mem[858] = 10'h370;
        mem[859] = 10'h02f;
        mem[860] = 10'h07b;
        mem[861] = 10'h3c0;
        mem[862] = 10'h36c;
        mem[863] = 10'h3d1;
        mem[864] = 10'h17b;
        mem[865] = 10'h388;
        mem[866] = 10'h32e;
        mem[867] = 10'h3ab;
        mem[868] = 10'h3cb;
        mem[869] = 10'h130;
        mem[870] = 10'h170;
        mem[871] = 10'h0c0;
        mem[872] = 10'h096;
        mem[873] = 10'h160;
        mem[874] = 10'h1e7;
        mem[875] = 10'h282;
        mem[876] = 10'h1f7;
        mem[877] = 10'h0de;
        mem[878] = 10'h106;
        mem[879] = 10'h184;
        mem[880] = 10'h081;
        mem[881] = 10'h3f7;
        mem[882] = 10'h373;
        mem[883] = 10'h1aa;
        mem[884] = 10'h380;
        mem[885] = 10'h14e;
        mem[886] = 10'h045;
        mem[887] = 10'h1eb;
        mem[888] = 10'h384;
        mem[889] = 10'h159;
        mem[890] = 10'h397;
        mem[891] = 10'h31e;
        mem[892] = 10'h0ba;
        mem[893] = 10'h1cd;
        mem[894] = 10'h3ef;
        mem[895] = 10'h0fa;
        mem[896] = 10'h06f;
        mem[897] = 10'h11d;
        mem[898] = 10'h233;
        mem[899] = 10'h287;
        mem[900] = 10'h235;
        mem[901] = 10'h049;
        mem[902] = 10'h2fc;
        mem[903] = 10'h39f;
        mem[904] = 10'h091;
        mem[905] = 10'h1d8;
        mem[906] = 10'h194;
        mem[907] = 10'h336;
        mem[908] = 10'h03d;
        mem[909] = 10'h1c1;
        mem[910] = 10'h2d5;
        mem[911] = 10'h2f8;
        mem[912] = 10'h14d;
        mem[913] = 10'h255;
        mem[914] = 10'h17f;
        mem[915] = 10'h245;
        mem[916] = 10'h219;
        mem[917] = 10'h0b7;
        mem[918] = 10'h2ab;
        mem[919] = 10'h01c;
        mem[920] = 10'h3ca;
        mem[921] = 10'h37a;
        mem[922] = 10'h1ef;
        mem[923] = 10'h231;
        mem[924] = 10'h3c4;
        mem[925] = 10'h2dd;
        mem[926] = 10'h039;
        mem[927] = 10'h1d6;
        mem[928] = 10'h1d1;
        mem[929] = 10'h0e6;
        mem[930] = 10'h263;
        mem[931] = 10'h190;
        mem[932] = 10'h0d7;
        mem[933] = 10'h0ca;
        mem[934] = 10'h23d;
        mem[935] = 10'h2de;
        mem[936] = 10'h1ad;
        mem[937] = 10'h36d;
        mem[938] = 10'h2ca;
        mem[939] = 10'h355;
        mem[940] = 10'h0ac;
        mem[941] = 10'h0db;
        mem[942] = 10'h128;
        mem[943] = 10'h0df;
        mem[944] = 10'h18f;
        mem[945] = 10'h3f2;
        mem[946] = 10'h037;
        mem[947] = 10'h115;
        mem[948] = 10'h35d;
        mem[949] = 10'h23b;
        mem[950] = 10'h1a6;
        mem[951] = 10'h2da;
        mem[952] = 10'h17a;
        mem[953] = 10'h1bb;
        mem[954] = 10'h0f9;
        mem[955] = 10'h28c;
        mem[956] = 10'h3dd;
        mem[957] = 10'h3f9;
        mem[958] = 10'h3a8;
        mem[959] = 10'h25f;
        mem[960] = 10'h07a;
        mem[961] = 10'h10c;
        mem[962] = 10'h120;
        mem[963] = 10'h090;
        mem[964] = 10'h0c1;
        mem[965] = 10'h047;
        mem[966] = 10'h15f;
        mem[967] = 10'h363;
        mem[968] = 10'h239;
        mem[969] = 10'h3a9;
        mem[970] = 10'h24c;
        mem[971] = 10'h31a;
        mem[972] = 10'h3c3;
        mem[973] = 10'h131;
        mem[974] = 10'h35a;
        mem[975] = 10'h0fd;
        mem[976] = 10'h172;
        mem[977] = 10'h3bc;
        mem[978] = 10'h18e;
        mem[979] = 10'h13e;
        mem[980] = 10'h142;
        mem[981] = 10'h22f;
        mem[982] = 10'h111;
        mem[983] = 10'h124;
        mem[984] = 10'h11e;
        mem[985] = 10'h1f4;
        mem[986] = 10'h11a;
        mem[987] = 10'h22c;
        mem[988] = 10'h3e4;
        mem[989] = 10'h009;
        mem[990] = 10'h372;
        mem[991] = 10'h157;
        mem[992] = 10'h382;
        mem[993] = 10'h0b1;
        mem[994] = 10'h3b4;
        mem[995] = 10'h242;
        mem[996] = 10'h2ad;
        mem[997] = 10'h3b1;
        mem[998] = 10'h261;
        mem[999] = 10'h112;
        mem[1000] = 10'h2c3;
        mem[1001] = 10'h312;
        mem[1002] = 10'h08a;
        mem[1003] = 10'h042;
        mem[1004] = 10'h34b;
        mem[1005] = 10'h0c9;
        mem[1006] = 10'h033;
        mem[1007] = 10'h25b;
        mem[1008] = 10'h046;
        mem[1009] = 10'h3e1;
        mem[1010] = 10'h0d5;
        mem[1011] = 10'h00a;
        mem[1012] = 10'h23e;
        mem[1013] = 10'h15a;
        mem[1014] = 10'h220;
        mem[1015] = 10'h1e0;
        mem[1016] = 10'h31f;
        mem[1017] = 10'h02b;
        mem[1018] = 10'h099;
        mem[1019] = 10'h186;
        mem[1020] = 10'h3bf;
        mem[1021] = 10'h3b3;
        mem[1022] = 10'h1da;
        mem[1023] = 10'h2ba;
    end
endmodule

module encrypt_4sbox_large3(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h0bf;
        mem[1] = 10'h0f0;
        mem[2] = 10'h0b4;
        mem[3] = 10'h2ce;
        mem[4] = 10'h00a;
        mem[5] = 10'h251;
        mem[6] = 10'h123;
        mem[7] = 10'h022;
        mem[8] = 10'h011;
        mem[9] = 10'h1e1;
        mem[10] = 10'h236;
        mem[11] = 10'h024;
        mem[12] = 10'h26b;
        mem[13] = 10'h322;
        mem[14] = 10'h025;
        mem[15] = 10'h13e;
        mem[16] = 10'h002;
        mem[17] = 10'h203;
        mem[18] = 10'h390;
        mem[19] = 10'h3bd;
        mem[20] = 10'h385;
        mem[21] = 10'h2db;
        mem[22] = 10'h069;
        mem[23] = 10'h25e;
        mem[24] = 10'h3a8;
        mem[25] = 10'h163;
        mem[26] = 10'h054;
        mem[27] = 10'h18d;
        mem[28] = 10'h3f8;
        mem[29] = 10'h18f;
        mem[30] = 10'h3f0;
        mem[31] = 10'h218;
        mem[32] = 10'h1c4;
        mem[33] = 10'h3a6;
        mem[34] = 10'h381;
        mem[35] = 10'h118;
        mem[36] = 10'h1df;
        mem[37] = 10'h3e1;
        mem[38] = 10'h334;
        mem[39] = 10'h341;
        mem[40] = 10'h13c;
        mem[41] = 10'h07f;
        mem[42] = 10'h043;
        mem[43] = 10'h10e;
        mem[44] = 10'h06f;
        mem[45] = 10'h3cd;
        mem[46] = 10'h3e7;
        mem[47] = 10'h3b7;
        mem[48] = 10'h188;
        mem[49] = 10'h295;
        mem[50] = 10'h121;
        mem[51] = 10'h04c;
        mem[52] = 10'h201;
        mem[53] = 10'h039;
        mem[54] = 10'h2b6;
        mem[55] = 10'h261;
        mem[56] = 10'h3ec;
        mem[57] = 10'h0c6;
        mem[58] = 10'h162;
        mem[59] = 10'h1e2;
        mem[60] = 10'h1ee;
        mem[61] = 10'h1ba;
        mem[62] = 10'h084;
        mem[63] = 10'h0a0;
        mem[64] = 10'h175;
        mem[65] = 10'h2b0;
        mem[66] = 10'h140;
        mem[67] = 10'h09f;
        mem[68] = 10'h19d;
        mem[69] = 10'h36a;
        mem[70] = 10'h12e;
        mem[71] = 10'h27d;
        mem[72] = 10'h2f6;
        mem[73] = 10'h2b7;
        mem[74] = 10'h26f;
        mem[75] = 10'h138;
        mem[76] = 10'h0c3;
        mem[77] = 10'h183;
        mem[78] = 10'h013;
        mem[79] = 10'h083;
        mem[80] = 10'h1f8;
        mem[81] = 10'h20f;
        mem[82] = 10'h3c3;
        mem[83] = 10'h184;
        mem[84] = 10'h030;
        mem[85] = 10'h1c5;
        mem[86] = 10'h0f6;
        mem[87] = 10'h03f;
        mem[88] = 10'h3ea;
        mem[89] = 10'h24f;
        mem[90] = 10'h009;
        mem[91] = 10'h231;
        mem[92] = 10'h2f8;
        mem[93] = 10'h016;
        mem[94] = 10'h181;
        mem[95] = 10'h30e;
        mem[96] = 10'h0c0;
        mem[97] = 10'h051;
        mem[98] = 10'h3fe;
        mem[99] = 10'h36c;
        mem[100] = 10'h1bb;
        mem[101] = 10'h370;
        mem[102] = 10'h290;
        mem[103] = 10'h098;
        mem[104] = 10'h303;
        mem[105] = 10'h03a;
        mem[106] = 10'h315;
        mem[107] = 10'h057;
        mem[108] = 10'h26d;
        mem[109] = 10'h22a;
        mem[110] = 10'h173;
        mem[111] = 10'h0ce;
        mem[112] = 10'h35f;
        mem[113] = 10'h226;
        mem[114] = 10'h1af;
        mem[115] = 10'h3ba;
        mem[116] = 10'h219;
        mem[117] = 10'h369;
        mem[118] = 10'h214;
        mem[119] = 10'h221;
        mem[120] = 10'h38e;
        mem[121] = 10'h2d9;
        mem[122] = 10'h29b;
        mem[123] = 10'h1f1;
        mem[124] = 10'h359;
        mem[125] = 10'h110;
        mem[126] = 10'h265;
        mem[127] = 10'h02a;
        mem[128] = 10'h21b;
        mem[129] = 10'h262;
        mem[130] = 10'h27e;
        mem[131] = 10'h1da;
        mem[132] = 10'h11d;
        mem[133] = 10'h159;
        mem[134] = 10'h092;
        mem[135] = 10'h08e;
        mem[136] = 10'h0e1;
        mem[137] = 10'h3c0;
        mem[138] = 10'h193;
        mem[139] = 10'h2b9;
        mem[140] = 10'h25d;
        mem[141] = 10'h353;
        mem[142] = 10'h033;
        mem[143] = 10'h350;
        mem[144] = 10'h367;
        mem[145] = 10'h0bb;
        mem[146] = 10'h310;
        mem[147] = 10'h23f;
        mem[148] = 10'h19c;
        mem[149] = 10'h260;
        mem[150] = 10'h1a7;
        mem[151] = 10'h151;
        mem[152] = 10'h332;
        mem[153] = 10'h142;
        mem[154] = 10'h052;
        mem[155] = 10'h1fe;
        mem[156] = 10'h2a2;
        mem[157] = 10'h2ab;
        mem[158] = 10'h16f;
        mem[159] = 10'h194;
        mem[160] = 10'h3d6;
        mem[161] = 10'h04a;
        mem[162] = 10'h23b;
        mem[163] = 10'h0d3;
        mem[164] = 10'h3d7;
        mem[165] = 10'h01d;
        mem[166] = 10'h13b;
        mem[167] = 10'h243;
        mem[168] = 10'h3a4;
        mem[169] = 10'h356;
        mem[170] = 10'h2b5;
        mem[171] = 10'h1e4;
        mem[172] = 10'h311;
        mem[173] = 10'h042;
        mem[174] = 10'h1f5;
        mem[175] = 10'h297;
        mem[176] = 10'h30b;
        mem[177] = 10'h1ec;
        mem[178] = 10'h39f;
        mem[179] = 10'h049;
        mem[180] = 10'h21e;
        mem[181] = 10'h22d;
        mem[182] = 10'h2bc;
        mem[183] = 10'h2fb;
        mem[184] = 10'h3a2;
        mem[185] = 10'h11b;
        mem[186] = 10'h132;
        mem[187] = 10'h333;
        mem[188] = 10'h16b;
        mem[189] = 10'h376;
        mem[190] = 10'h10d;
        mem[191] = 10'h28d;
        mem[192] = 10'h317;
        mem[193] = 10'h0b3;
        mem[194] = 10'h03b;
        mem[195] = 10'h1fc;
        mem[196] = 10'h2c0;
        mem[197] = 10'h2a6;
        mem[198] = 10'h143;
        mem[199] = 10'h0e9;
        mem[200] = 10'h3d4;
        mem[201] = 10'h055;
        mem[202] = 10'h32d;
        mem[203] = 10'h044;
        mem[204] = 10'h3c2;
        mem[205] = 10'h08d;
        mem[206] = 10'h0f5;
        mem[207] = 10'h16c;
        mem[208] = 10'h18e;
        mem[209] = 10'h2bf;
        mem[210] = 10'h18c;
        mem[211] = 10'h324;
        mem[212] = 10'h2a4;
        mem[213] = 10'h01e;
        mem[214] = 10'h102;
        mem[215] = 10'h1e3;
        mem[216] = 10'h02c;
        mem[217] = 10'h1d5;
        mem[218] = 10'h0d1;
        mem[219] = 10'h32e;
        mem[220] = 10'h010;
        mem[221] = 10'h0d8;
        mem[222] = 10'h0c7;
        mem[223] = 10'h3ef;
        mem[224] = 10'h22c;
        mem[225] = 10'h20c;
        mem[226] = 10'h397;
        mem[227] = 10'h050;
        mem[228] = 10'h0d9;
        mem[229] = 10'h33f;
        mem[230] = 10'h1c0;
        mem[231] = 10'h321;
        mem[232] = 10'h3c9;
        mem[233] = 10'h3a0;
        mem[234] = 10'h225;
        mem[235] = 10'h2ff;
        mem[236] = 10'h130;
        mem[237] = 10'h108;
        mem[238] = 10'h288;
        mem[239] = 10'h192;
        mem[240] = 10'h090;
        mem[241] = 10'h095;
        mem[242] = 10'h287;
        mem[243] = 10'h2be;
        mem[244] = 10'h1fa;
        mem[245] = 10'h0e5;
        mem[246] = 10'h0dc;
        mem[247] = 10'h32b;
        mem[248] = 10'h2c8;
        mem[249] = 10'h380;
        mem[250] = 10'h338;
        mem[251] = 10'h27f;
        mem[252] = 10'h3bc;
        mem[253] = 10'h314;
        mem[254] = 10'h3dc;
        mem[255] = 10'h1ab;
        mem[256] = 10'h388;
        mem[257] = 10'h25c;
        mem[258] = 10'h27c;
        mem[259] = 10'h1d2;
        mem[260] = 10'h1a4;
        mem[261] = 10'h1fd;
        mem[262] = 10'h339;
        mem[263] = 10'h294;
        mem[264] = 10'h389;
        mem[265] = 10'h23d;
        mem[266] = 10'h3a7;
        mem[267] = 10'h0e6;
        mem[268] = 10'h067;
        mem[269] = 10'h116;
        mem[270] = 10'h2f1;
        mem[271] = 10'h114;
        mem[272] = 10'h05f;
        mem[273] = 10'h0a3;
        mem[274] = 10'h1d7;
        mem[275] = 10'h377;
        mem[276] = 10'h36b;
        mem[277] = 10'h268;
        mem[278] = 10'h1ed;
        mem[279] = 10'h33a;
        mem[280] = 10'h1c3;
        mem[281] = 10'h2dd;
        mem[282] = 10'h3de;
        mem[283] = 10'h379;
        mem[284] = 10'h139;
        mem[285] = 10'h305;
        mem[286] = 10'h22e;
        mem[287] = 10'h3e4;
        mem[288] = 10'h08c;
        mem[289] = 10'h007;
        mem[290] = 10'h363;
        mem[291] = 10'h004;
        mem[292] = 10'h185;
        mem[293] = 10'h255;
        mem[294] = 10'h365;
        mem[295] = 10'h357;
        mem[296] = 10'h2fd;
        mem[297] = 10'h2c4;
        mem[298] = 10'h38b;
        mem[299] = 10'h0a2;
        mem[300] = 10'h106;
        mem[301] = 10'h3cc;
        mem[302] = 10'h0aa;
        mem[303] = 10'h3e9;
        mem[304] = 10'h202;
        mem[305] = 10'h271;
        mem[306] = 10'h019;
        mem[307] = 10'h26e;
        mem[308] = 10'h344;
        mem[309] = 10'h331;
        mem[310] = 10'h1b9;
        mem[311] = 10'h2bb;
        mem[312] = 10'h313;
        mem[313] = 10'h2e1;
        mem[314] = 10'h1d3;
        mem[315] = 10'h1b0;
        mem[316] = 10'h3d1;
        mem[317] = 10'h386;
        mem[318] = 10'h27a;
        mem[319] = 10'h3ce;
        mem[320] = 10'h0d5;
        mem[321] = 10'h3c7;
        mem[322] = 10'h087;
        mem[323] = 10'h235;
        mem[324] = 10'h14b;
        mem[325] = 10'h269;
        mem[326] = 10'h25f;
        mem[327] = 10'h2f0;
        mem[328] = 10'h047;
        mem[329] = 10'h2fe;
        mem[330] = 10'h299;
        mem[331] = 10'h197;
        mem[332] = 10'h34c;
        mem[333] = 10'h003;
        mem[334] = 10'h0ae;
        mem[335] = 10'h39d;
        mem[336] = 10'h335;
        mem[337] = 10'h0ec;
        mem[338] = 10'h01c;
        mem[339] = 10'h2ae;
        mem[340] = 10'h1e5;
        mem[341] = 10'h15f;
        mem[342] = 10'h1c8;
        mem[343] = 10'h06d;
        mem[344] = 10'h2f2;
        mem[345] = 10'h2d5;
        mem[346] = 10'h17b;
        mem[347] = 10'h3e2;
        mem[348] = 10'h228;
        mem[349] = 10'h1eb;
        mem[350] = 10'h0cc;
        mem[351] = 10'h147;
        mem[352] = 10'h00b;
        mem[353] = 10'h3f1;
        mem[354] = 10'h125;
        mem[355] = 10'h20e;
        mem[356] = 10'h0ef;
        mem[357] = 10'h21a;
        mem[358] = 10'h0b7;
        mem[359] = 10'h204;
        mem[360] = 10'h2cc;
        mem[361] = 10'h3f6;
        mem[362] = 10'h1ce;
        mem[363] = 10'h031;
        mem[364] = 10'h0fa;
        mem[365] = 10'h127;
        mem[366] = 10'h152;
        mem[367] = 10'h064;
        mem[368] = 10'h358;
        mem[369] = 10'h086;
        mem[370] = 10'h3eb;
        mem[371] = 10'h222;
        mem[372] = 10'h20a;
        mem[373] = 10'h2af;
        mem[374] = 10'h325;
        mem[375] = 10'h2cb;
        mem[376] = 10'h01b;
        mem[377] = 10'h072;
        mem[378] = 10'h11f;
        mem[379] = 10'h00d;
        mem[380] = 10'h336;
        mem[381] = 10'h3c8;
        mem[382] = 10'h31b;
        mem[383] = 10'h2e7;
        mem[384] = 10'h282;
        mem[385] = 10'h060;
        mem[386] = 10'h1f6;
        mem[387] = 10'h32a;
        mem[388] = 10'h158;
        mem[389] = 10'h39b;
        mem[390] = 10'h0dd;
        mem[391] = 10'h323;
        mem[392] = 10'h3e0;
        mem[393] = 10'h3ca;
        mem[394] = 10'h22b;
        mem[395] = 10'h238;
        mem[396] = 10'h10b;
        mem[397] = 10'h246;
        mem[398] = 10'h3c6;
        mem[399] = 10'h35d;
        mem[400] = 10'h29e;
        mem[401] = 10'h32f;
        mem[402] = 10'h0e2;
        mem[403] = 10'h29d;
        mem[404] = 10'h063;
        mem[405] = 10'h368;
        mem[406] = 10'h382;
        mem[407] = 10'h15a;
        mem[408] = 10'h2a0;
        mem[409] = 10'h0e8;
        mem[410] = 10'h18a;
        mem[411] = 10'h176;
        mem[412] = 10'h318;
        mem[413] = 10'h15b;
        mem[414] = 10'h0cf;
        mem[415] = 10'h06c;
        mem[416] = 10'h145;
        mem[417] = 10'h3c4;
        mem[418] = 10'h351;
        mem[419] = 10'h1fb;
        mem[420] = 10'h1dc;
        mem[421] = 10'h259;
        mem[422] = 10'h1d0;
        mem[423] = 10'h373;
        mem[424] = 10'h0e3;
        mem[425] = 10'h1c7;
        mem[426] = 10'h240;
        mem[427] = 10'h31c;
        mem[428] = 10'h33d;
        mem[429] = 10'h093;
        mem[430] = 10'h36f;
        mem[431] = 10'h2d3;
        mem[432] = 10'h0ab;
        mem[433] = 10'h05d;
        mem[434] = 10'h029;
        mem[435] = 10'h34f;
        mem[436] = 10'h00c;
        mem[437] = 10'h31f;
        mem[438] = 10'h38c;
        mem[439] = 10'h2dc;
        mem[440] = 10'h26c;
        mem[441] = 10'h1e7;
        mem[442] = 10'h34a;
        mem[443] = 10'h29c;
        mem[444] = 10'h070;
        mem[445] = 10'h12b;
        mem[446] = 10'h1bc;
        mem[447] = 10'h1a2;
        mem[448] = 10'h0bc;
        mem[449] = 10'h12d;
        mem[450] = 10'h0ea;
        mem[451] = 10'h02f;
        mem[452] = 10'h347;
        mem[453] = 10'h2e3;
        mem[454] = 10'h250;
        mem[455] = 10'h2eb;
        mem[456] = 10'h0f3;
        mem[457] = 10'h062;
        mem[458] = 10'h39e;
        mem[459] = 10'h02d;
        mem[460] = 10'h015;
        mem[461] = 10'h14e;
        mem[462] = 10'h2de;
        mem[463] = 10'h1a8;
        mem[464] = 10'h1f4;
        mem[465] = 10'h247;
        mem[466] = 10'h099;
        mem[467] = 10'h014;
        mem[468] = 10'h0d4;
        mem[469] = 10'h2d6;
        mem[470] = 10'h1ae;
        mem[471] = 10'h191;
        mem[472] = 10'h3c5;
        mem[473] = 10'h208;
        mem[474] = 10'h2e0;
        mem[475] = 10'h01f;
        mem[476] = 10'h2c7;
        mem[477] = 10'h25b;
        mem[478] = 10'h171;
        mem[479] = 10'h2b3;
        mem[480] = 10'h1db;
        mem[481] = 10'h195;
        mem[482] = 10'h122;
        mem[483] = 10'h2d8;
        mem[484] = 10'h2ac;
        mem[485] = 10'h0a1;
        mem[486] = 10'h2ba;
        mem[487] = 10'h0b2;
        mem[488] = 10'h337;
        mem[489] = 10'h144;
        mem[490] = 10'h252;
        mem[491] = 10'h021;
        mem[492] = 10'h131;
        mem[493] = 10'h309;
        mem[494] = 10'h26a;
        mem[495] = 10'h06e;
        mem[496] = 10'h326;
        mem[497] = 10'h304;
        mem[498] = 10'h2a1;
        mem[499] = 10'h360;
        mem[500] = 10'h0f4;
        mem[501] = 10'h398;
        mem[502] = 10'h229;
        mem[503] = 10'h237;
        mem[504] = 10'h115;
        mem[505] = 10'h37f;
        mem[506] = 10'h234;
        mem[507] = 10'h38a;
        mem[508] = 10'h2e2;
        mem[509] = 10'h153;
        mem[510] = 10'h232;
        mem[511] = 10'h089;
        mem[512] = 10'h187;
        mem[513] = 10'h1a9;
        mem[514] = 10'h0db;
        mem[515] = 10'h136;
        mem[516] = 10'h2c1;
        mem[517] = 10'h2ed;
        mem[518] = 10'h11e;
        mem[519] = 10'h071;
        mem[520] = 10'h1ca;
        mem[521] = 10'h2a5;
        mem[522] = 10'h161;
        mem[523] = 10'h0a9;
        mem[524] = 10'h0b8;
        mem[525] = 10'h3bf;
        mem[526] = 10'h1b6;
        mem[527] = 10'h05c;
        mem[528] = 10'h07b;
        mem[529] = 10'h300;
        mem[530] = 10'h3fa;
        mem[531] = 10'h155;
        mem[532] = 10'h3f5;
        mem[533] = 10'h316;
        mem[534] = 10'h046;
        mem[535] = 10'h034;
        mem[536] = 10'h2d4;
        mem[537] = 10'h074;
        mem[538] = 10'h263;
        mem[539] = 10'h1a1;
        mem[540] = 10'h24b;
        mem[541] = 10'h307;
        mem[542] = 10'h1bd;
        mem[543] = 10'h0ff;
        mem[544] = 10'h023;
        mem[545] = 10'h008;
        mem[546] = 10'h3b1;
        mem[547] = 10'h05a;
        mem[548] = 10'h053;
        mem[549] = 10'h340;
        mem[550] = 10'h124;
        mem[551] = 10'h3e5;
        mem[552] = 10'h3b9;
        mem[553] = 10'h09e;
        mem[554] = 10'h17d;
        mem[555] = 10'h1c6;
        mem[556] = 10'h270;
        mem[557] = 10'h1ac;
        mem[558] = 10'h1ea;
        mem[559] = 10'h366;
        mem[560] = 10'h006;
        mem[561] = 10'h1aa;
        mem[562] = 10'h0fd;
        mem[563] = 10'h283;
        mem[564] = 10'h0cd;
        mem[565] = 10'h20d;
        mem[566] = 10'h29a;
        mem[567] = 10'h217;
        mem[568] = 10'h129;
        mem[569] = 10'h0ed;
        mem[570] = 10'h18b;
        mem[571] = 10'h168;
        mem[572] = 10'h371;
        mem[573] = 10'h1e9;
        mem[574] = 10'h2d7;
        mem[575] = 10'h391;
        mem[576] = 10'h04d;
        mem[577] = 10'h230;
        mem[578] = 10'h3d5;
        mem[579] = 10'h39c;
        mem[580] = 10'h2f3;
        mem[581] = 10'h0f2;
        mem[582] = 10'h3c1;
        mem[583] = 10'h076;
        mem[584] = 10'h2ca;
        mem[585] = 10'h35c;
        mem[586] = 10'h2ec;
        mem[587] = 10'h206;
        mem[588] = 10'h05b;
        mem[589] = 10'h296;
        mem[590] = 10'h0eb;
        mem[591] = 10'h16d;
        mem[592] = 10'h36d;
        mem[593] = 10'h0b0;
        mem[594] = 10'h11c;
        mem[595] = 10'h3ff;
        mem[596] = 10'h2ee;
        mem[597] = 10'h03e;
        mem[598] = 10'h308;
        mem[599] = 10'h2a7;
        mem[600] = 10'h134;
        mem[601] = 10'h0fe;
        mem[602] = 10'h20b;
        mem[603] = 10'h3ad;
        mem[604] = 10'h1a6;
        mem[605] = 10'h040;
        mem[606] = 10'h3d8;
        mem[607] = 10'h343;
        mem[608] = 10'h276;
        mem[609] = 10'h0a4;
        mem[610] = 10'h2da;
        mem[611] = 10'h2cf;
        mem[612] = 10'h0be;
        mem[613] = 10'h177;
        mem[614] = 10'h1cd;
        mem[615] = 10'h1b5;
        mem[616] = 10'h005;
        mem[617] = 10'h23a;
        mem[618] = 10'h048;
        mem[619] = 10'h2f5;
        mem[620] = 10'h1a5;
        mem[621] = 10'h2f7;
        mem[622] = 10'h223;
        mem[623] = 10'h256;
        mem[624] = 10'h028;
        mem[625] = 10'h09a;
        mem[626] = 10'h0af;
        mem[627] = 10'h2f4;
        mem[628] = 10'h2ea;
        mem[629] = 10'h3b2;
        mem[630] = 10'h2b1;
        mem[631] = 10'h2c6;
        mem[632] = 10'h327;
        mem[633] = 10'h1d1;
        mem[634] = 10'h1f9;
        mem[635] = 10'h1f2;
        mem[636] = 10'h205;
        mem[637] = 10'h3a5;
        mem[638] = 10'h07c;
        mem[639] = 10'h281;
        mem[640] = 10'h399;
        mem[641] = 10'h180;
        mem[642] = 10'h241;
        mem[643] = 10'h198;
        mem[644] = 10'h104;
        mem[645] = 10'h094;
        mem[646] = 10'h0d6;
        mem[647] = 10'h3b3;
        mem[648] = 10'h2b4;
        mem[649] = 10'h02b;
        mem[650] = 10'h372;
        mem[651] = 10'h169;
        mem[652] = 10'h3ae;
        mem[653] = 10'h133;
        mem[654] = 10'h1d6;
        mem[655] = 10'h2e4;
        mem[656] = 10'h065;
        mem[657] = 10'h37a;
        mem[658] = 10'h37c;
        mem[659] = 10'h08b;
        mem[660] = 10'h036;
        mem[661] = 10'h2d2;
        mem[662] = 10'h17c;
        mem[663] = 10'h150;
        mem[664] = 10'h375;
        mem[665] = 10'h3d0;
        mem[666] = 10'h0b9;
        mem[667] = 10'h1b8;
        mem[668] = 10'h254;
        mem[669] = 10'h19e;
        mem[670] = 10'h2b8;
        mem[671] = 10'h166;
        mem[672] = 10'h289;
        mem[673] = 10'h13f;
        mem[674] = 10'h160;
        mem[675] = 10'h15c;
        mem[676] = 10'h04b;
        mem[677] = 10'h3f9;
        mem[678] = 10'h14d;
        mem[679] = 10'h33e;
        mem[680] = 10'h2d1;
        mem[681] = 10'h012;
        mem[682] = 10'h330;
        mem[683] = 10'h0e0;
        mem[684] = 10'h038;
        mem[685] = 10'h36e;
        mem[686] = 10'h026;
        mem[687] = 10'h1d8;
        mem[688] = 10'h045;
        mem[689] = 10'h2c9;
        mem[690] = 10'h027;
        mem[691] = 10'h392;
        mem[692] = 10'h146;
        mem[693] = 10'h1a3;
        mem[694] = 10'h2e6;
        mem[695] = 10'h135;
        mem[696] = 10'h25a;
        mem[697] = 10'h2f9;
        mem[698] = 10'h0b5;
        mem[699] = 10'h2ad;
        mem[700] = 10'h126;
        mem[701] = 10'h16a;
        mem[702] = 10'h384;
        mem[703] = 10'h1ef;
        mem[704] = 10'h182;
        mem[705] = 10'h396;
        mem[706] = 10'h1d4;
        mem[707] = 10'h109;
        mem[708] = 10'h19b;
        mem[709] = 10'h30c;
        mem[710] = 10'h3d2;
        mem[711] = 10'h2a3;
        mem[712] = 10'h1ff;
        mem[713] = 10'h274;
        mem[714] = 10'h149;
        mem[715] = 10'h286;
        mem[716] = 10'h2a9;
        mem[717] = 10'h3f4;
        mem[718] = 10'h2c2;
        mem[719] = 10'h13d;
        mem[720] = 10'h167;
        mem[721] = 10'h2b2;
        mem[722] = 10'h362;
        mem[723] = 10'h15e;
        mem[724] = 10'h38d;
        mem[725] = 10'h186;
        mem[726] = 10'h0f9;
        mem[727] = 10'h3e8;
        mem[728] = 10'h301;
        mem[729] = 10'h2e8;
        mem[730] = 10'h292;
        mem[731] = 10'h345;
        mem[732] = 10'h03c;
        mem[733] = 10'h3ee;
        mem[734] = 10'h157;
        mem[735] = 10'h080;
        mem[736] = 10'h032;
        mem[737] = 10'h1e6;
        mem[738] = 10'h085;
        mem[739] = 10'h3d9;
        mem[740] = 10'h3f2;
        mem[741] = 10'h00e;
        mem[742] = 10'h0fb;
        mem[743] = 10'h101;
        mem[744] = 10'h1c1;
        mem[745] = 10'h249;
        mem[746] = 10'h39a;
        mem[747] = 10'h00f;
        mem[748] = 10'h128;
        mem[749] = 10'h07d;
        mem[750] = 10'h10a;
        mem[751] = 10'h209;
        mem[752] = 10'h329;
        mem[753] = 10'h393;
        mem[754] = 10'h2c3;
        mem[755] = 10'h2d0;
        mem[756] = 10'h097;
        mem[757] = 10'h34e;
        mem[758] = 10'h05e;
        mem[759] = 10'h30f;
        mem[760] = 10'h266;
        mem[761] = 10'h0d0;
        mem[762] = 10'h1cf;
        mem[763] = 10'h28e;
        mem[764] = 10'h28b;
        mem[765] = 10'h37d;
        mem[766] = 10'h107;
        mem[767] = 10'h078;
        mem[768] = 10'h24a;
        mem[769] = 10'h091;
        mem[770] = 10'h0df;
        mem[771] = 10'h1d9;
        mem[772] = 10'h3fc;
        mem[773] = 10'h1e0;
        mem[774] = 10'h346;
        mem[775] = 10'h253;
        mem[776] = 10'h0ee;
        mem[777] = 10'h24d;
        mem[778] = 10'h0b6;
        mem[779] = 10'h21d;
        mem[780] = 10'h08a;
        mem[781] = 10'h1b1;
        mem[782] = 10'h302;
        mem[783] = 10'h1de;
        mem[784] = 10'h079;
        mem[785] = 10'h07a;
        mem[786] = 10'h3be;
        mem[787] = 10'h3e3;
        mem[788] = 10'h1e8;
        mem[789] = 10'h0ad;
        mem[790] = 10'h3f3;
        mem[791] = 10'h1f7;
        mem[792] = 10'h117;
        mem[793] = 10'h081;
        mem[794] = 10'h15d;
        mem[795] = 10'h273;
        mem[796] = 10'h216;
        mem[797] = 10'h3da;
        mem[798] = 10'h23e;
        mem[799] = 10'h27b;
        mem[800] = 10'h1f0;
        mem[801] = 10'h112;
        mem[802] = 10'h09c;
        mem[803] = 10'h16e;
        mem[804] = 10'h001;
        mem[805] = 10'h3e6;
        mem[806] = 10'h320;
        mem[807] = 10'h0a7;
        mem[808] = 10'h242;
        mem[809] = 10'h34d;
        mem[810] = 10'h189;
        mem[811] = 10'h0c9;
        mem[812] = 10'h28a;
        mem[813] = 10'h395;
        mem[814] = 10'h2cd;
        mem[815] = 10'h196;
        mem[816] = 10'h020;
        mem[817] = 10'h224;
        mem[818] = 10'h0d7;
        mem[819] = 10'h348;
        mem[820] = 10'h342;
        mem[821] = 10'h28f;
        mem[822] = 10'h165;
        mem[823] = 10'h3af;
        mem[824] = 10'h239;
        mem[825] = 10'h3b4;
        mem[826] = 10'h035;
        mem[827] = 10'h258;
        mem[828] = 10'h21f;
        mem[829] = 10'h075;
        mem[830] = 10'h30a;
        mem[831] = 10'h200;
        mem[832] = 10'h2fc;
        mem[833] = 10'h14a;
        mem[834] = 10'h3b5;
        mem[835] = 10'h14c;
        mem[836] = 10'h018;
        mem[837] = 10'h1cb;
        mem[838] = 10'h1be;
        mem[839] = 10'h2e9;
        mem[840] = 10'h0bd;
        mem[841] = 10'h0d2;
        mem[842] = 10'h148;
        mem[843] = 10'h10f;
        mem[844] = 10'h1ad;
        mem[845] = 10'h0c5;
        mem[846] = 10'h0e4;
        mem[847] = 10'h3df;
        mem[848] = 10'h3dd;
        mem[849] = 10'h17e;
        mem[850] = 10'h061;
        mem[851] = 10'h257;
        mem[852] = 10'h3a3;
        mem[853] = 10'h244;
        mem[854] = 10'h3ed;
        mem[855] = 10'h37b;
        mem[856] = 10'h32c;
        mem[857] = 10'h10c;
        mem[858] = 10'h23c;
        mem[859] = 10'h3b6;
        mem[860] = 10'h082;
        mem[861] = 10'h0ba;
        mem[862] = 10'h227;
        mem[863] = 10'h211;
        mem[864] = 10'h164;
        mem[865] = 10'h279;
        mem[866] = 10'h213;
        mem[867] = 10'h293;
        mem[868] = 10'h172;
        mem[869] = 10'h215;
        mem[870] = 10'h190;
        mem[871] = 10'h105;
        mem[872] = 10'h245;
        mem[873] = 10'h04e;
        mem[874] = 10'h33c;
        mem[875] = 10'h12c;
        mem[876] = 10'h387;
        mem[877] = 10'h291;
        mem[878] = 10'h349;
        mem[879] = 10'h037;
        mem[880] = 10'h06b;
        mem[881] = 10'h000;
        mem[882] = 10'h394;
        mem[883] = 10'h22f;
        mem[884] = 10'h3aa;
        mem[885] = 10'h17f;
        mem[886] = 10'h179;
        mem[887] = 10'h31e;
        mem[888] = 10'h28c;
        mem[889] = 10'h0ca;
        mem[890] = 10'h0c2;
        mem[891] = 10'h077;
        mem[892] = 10'h319;
        mem[893] = 10'h14f;
        mem[894] = 10'h2e5;
        mem[895] = 10'h37e;
        mem[896] = 10'h073;
        mem[897] = 10'h3bb;
        mem[898] = 10'h298;
        mem[899] = 10'h0fc;
        mem[900] = 10'h2aa;
        mem[901] = 10'h3f7;
        mem[902] = 10'h120;
        mem[903] = 10'h19f;
        mem[904] = 10'h1cc;
        mem[905] = 10'h1b2;
        mem[906] = 10'h2c5;
        mem[907] = 10'h30d;
        mem[908] = 10'h01a;
        mem[909] = 10'h0c1;
        mem[910] = 10'h17a;
        mem[911] = 10'h02e;
        mem[912] = 10'h354;
        mem[913] = 10'h1b3;
        mem[914] = 10'h154;
        mem[915] = 10'h1c2;
        mem[916] = 10'h0e7;
        mem[917] = 10'h156;
        mem[918] = 10'h3a1;
        mem[919] = 10'h0a8;
        mem[920] = 10'h119;
        mem[921] = 10'h3a9;
        mem[922] = 10'h017;
        mem[923] = 10'h0a5;
        mem[924] = 10'h264;
        mem[925] = 10'h355;
        mem[926] = 10'h056;
        mem[927] = 10'h284;
        mem[928] = 10'h0f8;
        mem[929] = 10'h113;
        mem[930] = 10'h220;
        mem[931] = 10'h3b0;
        mem[932] = 10'h12f;
        mem[933] = 10'h3ac;
        mem[934] = 10'h3fb;
        mem[935] = 10'h3db;
        mem[936] = 10'h066;
        mem[937] = 10'h04f;
        mem[938] = 10'h35e;
        mem[939] = 10'h31d;
        mem[940] = 10'h0f1;
        mem[941] = 10'h285;
        mem[942] = 10'h0f7;
        mem[943] = 10'h178;
        mem[944] = 10'h275;
        mem[945] = 10'h0c8;
        mem[946] = 10'h058;
        mem[947] = 10'h207;
        mem[948] = 10'h0de;
        mem[949] = 10'h378;
        mem[950] = 10'h07e;
        mem[951] = 10'h24c;
        mem[952] = 10'h088;
        mem[953] = 10'h3cb;
        mem[954] = 10'h103;
        mem[955] = 10'h03d;
        mem[956] = 10'h38f;
        mem[957] = 10'h2a8;
        mem[958] = 10'h352;
        mem[959] = 10'h137;
        mem[960] = 10'h3ab;
        mem[961] = 10'h212;
        mem[962] = 10'h13a;
        mem[963] = 10'h2ef;
        mem[964] = 10'h364;
        mem[965] = 10'h2df;
        mem[966] = 10'h233;
        mem[967] = 10'h267;
        mem[968] = 10'h111;
        mem[969] = 10'h3d3;
        mem[970] = 10'h1f3;
        mem[971] = 10'h1dd;
        mem[972] = 10'h361;
        mem[973] = 10'h278;
        mem[974] = 10'h100;
        mem[975] = 10'h1b7;
        mem[976] = 10'h2bd;
        mem[977] = 10'h280;
        mem[978] = 10'h0da;
        mem[979] = 10'h06a;
        mem[980] = 10'h141;
        mem[981] = 10'h374;
        mem[982] = 10'h08f;
        mem[983] = 10'h21c;
        mem[984] = 10'h12a;
        mem[985] = 10'h096;
        mem[986] = 10'h11a;
        mem[987] = 10'h383;
        mem[988] = 10'h0a6;
        mem[989] = 10'h09d;
        mem[990] = 10'h31a;
        mem[991] = 10'h35b;
        mem[992] = 10'h306;
        mem[993] = 10'h0c4;
        mem[994] = 10'h328;
        mem[995] = 10'h210;
        mem[996] = 10'h041;
        mem[997] = 10'h272;
        mem[998] = 10'h0cb;
        mem[999] = 10'h174;
        mem[1000] = 10'h1a0;
        mem[1001] = 10'h170;
        mem[1002] = 10'h3fd;
        mem[1003] = 10'h1b4;
        mem[1004] = 10'h312;
        mem[1005] = 10'h0ac;
        mem[1006] = 10'h1bf;
        mem[1007] = 10'h1c9;
        mem[1008] = 10'h3cf;
        mem[1009] = 10'h09b;
        mem[1010] = 10'h24e;
        mem[1011] = 10'h248;
        mem[1012] = 10'h29f;
        mem[1013] = 10'h19a;
        mem[1014] = 10'h199;
        mem[1015] = 10'h068;
        mem[1016] = 10'h2fa;
        mem[1017] = 10'h0b1;
        mem[1018] = 10'h3b8;
        mem[1019] = 10'h277;
        mem[1020] = 10'h33b;
        mem[1021] = 10'h35a;
        mem[1022] = 10'h059;
        mem[1023] = 10'h34b;
    end
endmodule

module encrypt_4sbox_large4(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h302;
        mem[1] = 10'h246;
        mem[2] = 10'h2f9;
        mem[3] = 10'h075;
        mem[4] = 10'h346;
        mem[5] = 10'h277;
        mem[6] = 10'h0c8;
        mem[7] = 10'h099;
        mem[8] = 10'h2f7;
        mem[9] = 10'h01e;
        mem[10] = 10'h128;
        mem[11] = 10'h08a;
        mem[12] = 10'h110;
        mem[13] = 10'h3f5;
        mem[14] = 10'h31f;
        mem[15] = 10'h1b8;
        mem[16] = 10'h03d;
        mem[17] = 10'h244;
        mem[18] = 10'h0b3;
        mem[19] = 10'h2d3;
        mem[20] = 10'h02b;
        mem[21] = 10'h23a;
        mem[22] = 10'h313;
        mem[23] = 10'h197;
        mem[24] = 10'h09e;
        mem[25] = 10'h129;
        mem[26] = 10'h216;
        mem[27] = 10'h0ef;
        mem[28] = 10'h3ee;
        mem[29] = 10'h2b6;
        mem[30] = 10'h34a;
        mem[31] = 10'h252;
        mem[32] = 10'h04b;
        mem[33] = 10'h2c5;
        mem[34] = 10'h1ef;
        mem[35] = 10'h1bb;
        mem[36] = 10'h27d;
        mem[37] = 10'h04d;
        mem[38] = 10'h054;
        mem[39] = 10'h3db;
        mem[40] = 10'h040;
        mem[41] = 10'h3d0;
        mem[42] = 10'h13e;
        mem[43] = 10'h2ce;
        mem[44] = 10'h2f1;
        mem[45] = 10'h2da;
        mem[46] = 10'h0fb;
        mem[47] = 10'h31a;
        mem[48] = 10'h278;
        mem[49] = 10'h06f;
        mem[50] = 10'h3ac;
        mem[51] = 10'h37a;
        mem[52] = 10'h074;
        mem[53] = 10'h135;
        mem[54] = 10'h35e;
        mem[55] = 10'h032;
        mem[56] = 10'h085;
        mem[57] = 10'h07b;
        mem[58] = 10'h303;
        mem[59] = 10'h207;
        mem[60] = 10'h38d;
        mem[61] = 10'h0d3;
        mem[62] = 10'h00e;
        mem[63] = 10'h298;
        mem[64] = 10'h316;
        mem[65] = 10'h0c3;
        mem[66] = 10'h213;
        mem[67] = 10'h01f;
        mem[68] = 10'h3d2;
        mem[69] = 10'h3e2;
        mem[70] = 10'h250;
        mem[71] = 10'h1b5;
        mem[72] = 10'h372;
        mem[73] = 10'h090;
        mem[74] = 10'h383;
        mem[75] = 10'h39b;
        mem[76] = 10'h0f0;
        mem[77] = 10'h023;
        mem[78] = 10'h376;
        mem[79] = 10'h0a0;
        mem[80] = 10'h157;
        mem[81] = 10'h1ab;
        mem[82] = 10'h1a1;
        mem[83] = 10'h035;
        mem[84] = 10'h194;
        mem[85] = 10'h04e;
        mem[86] = 10'h380;
        mem[87] = 10'h06e;
        mem[88] = 10'h367;
        mem[89] = 10'h274;
        mem[90] = 10'h186;
        mem[91] = 10'h314;
        mem[92] = 10'h10f;
        mem[93] = 10'h293;
        mem[94] = 10'h3fa;
        mem[95] = 10'h220;
        mem[96] = 10'h3b2;
        mem[97] = 10'h20b;
        mem[98] = 10'h15a;
        mem[99] = 10'h3b0;
        mem[100] = 10'h212;
        mem[101] = 10'h0a6;
        mem[102] = 10'h3a9;
        mem[103] = 10'h1be;
        mem[104] = 10'h13f;
        mem[105] = 10'h23b;
        mem[106] = 10'h3da;
        mem[107] = 10'h24e;
        mem[108] = 10'h113;
        mem[109] = 10'h38f;
        mem[110] = 10'h11e;
        mem[111] = 10'h00a;
        mem[112] = 10'h3af;
        mem[113] = 10'h236;
        mem[114] = 10'h368;
        mem[115] = 10'h15d;
        mem[116] = 10'h25e;
        mem[117] = 10'h317;
        mem[118] = 10'h149;
        mem[119] = 10'h12a;
        mem[120] = 10'h1dd;
        mem[121] = 10'h264;
        mem[122] = 10'h0ad;
        mem[123] = 10'h282;
        mem[124] = 10'h12e;
        mem[125] = 10'h139;
        mem[126] = 10'h05b;
        mem[127] = 10'h1d9;
        mem[128] = 10'h1e4;
        mem[129] = 10'h1e6;
        mem[130] = 10'h0eb;
        mem[131] = 10'h3df;
        mem[132] = 10'h0c1;
        mem[133] = 10'h358;
        mem[134] = 10'h12c;
        mem[135] = 10'h063;
        mem[136] = 10'h3a8;
        mem[137] = 10'h1a0;
        mem[138] = 10'h20a;
        mem[139] = 10'h161;
        mem[140] = 10'h001;
        mem[141] = 10'h2ef;
        mem[142] = 10'h3b4;
        mem[143] = 10'h17c;
        mem[144] = 10'h227;
        mem[145] = 10'h120;
        mem[146] = 10'h3a7;
        mem[147] = 10'h0a3;
        mem[148] = 10'h29b;
        mem[149] = 10'h0df;
        mem[150] = 10'h222;
        mem[151] = 10'h34c;
        mem[152] = 10'h1ee;
        mem[153] = 10'h053;
        mem[154] = 10'h33a;
        mem[155] = 10'h147;
        mem[156] = 10'h13b;
        mem[157] = 10'h200;
        mem[158] = 10'h153;
        mem[159] = 10'h0ca;
        mem[160] = 10'h337;
        mem[161] = 10'h1db;
        mem[162] = 10'h051;
        mem[163] = 10'h1ad;
        mem[164] = 10'h104;
        mem[165] = 10'h079;
        mem[166] = 10'h39f;
        mem[167] = 10'h14e;
        mem[168] = 10'h125;
        mem[169] = 10'h290;
        mem[170] = 10'h22a;
        mem[171] = 10'h0f6;
        mem[172] = 10'h1bf;
        mem[173] = 10'h272;
        mem[174] = 10'h2d5;
        mem[175] = 10'h3cf;
        mem[176] = 10'h036;
        mem[177] = 10'h029;
        mem[178] = 10'h05c;
        mem[179] = 10'h1d8;
        mem[180] = 10'h10b;
        mem[181] = 10'h1f6;
        mem[182] = 10'h185;
        mem[183] = 10'h078;
        mem[184] = 10'h191;
        mem[185] = 10'h3be;
        mem[186] = 10'h1d3;
        mem[187] = 10'h073;
        mem[188] = 10'h28e;
        mem[189] = 10'h08c;
        mem[190] = 10'h20f;
        mem[191] = 10'h390;
        mem[192] = 10'h25a;
        mem[193] = 10'h095;
        mem[194] = 10'h112;
        mem[195] = 10'h1b6;
        mem[196] = 10'h21e;
        mem[197] = 10'h031;
        mem[198] = 10'h177;
        mem[199] = 10'h2b7;
        mem[200] = 10'h3e4;
        mem[201] = 10'h32e;
        mem[202] = 10'h37c;
        mem[203] = 10'h26a;
        mem[204] = 10'h2fb;
        mem[205] = 10'h072;
        mem[206] = 10'h04c;
        mem[207] = 10'h36a;
        mem[208] = 10'h170;
        mem[209] = 10'h0ed;
        mem[210] = 10'h06c;
        mem[211] = 10'h357;
        mem[212] = 10'h06b;
        mem[213] = 10'h0e4;
        mem[214] = 10'h3c7;
        mem[215] = 10'h285;
        mem[216] = 10'h3d4;
        mem[217] = 10'h2ac;
        mem[218] = 10'h39c;
        mem[219] = 10'h311;
        mem[220] = 10'h2dc;
        mem[221] = 10'h101;
        mem[222] = 10'h219;
        mem[223] = 10'h152;
        mem[224] = 10'h3eb;
        mem[225] = 10'h2cf;
        mem[226] = 10'h27b;
        mem[227] = 10'h3ff;
        mem[228] = 10'h137;
        mem[229] = 10'h0e0;
        mem[230] = 10'h2ec;
        mem[231] = 10'h2ee;
        mem[232] = 10'h020;
        mem[233] = 10'h241;
        mem[234] = 10'h2fc;
        mem[235] = 10'h046;
        mem[236] = 10'h0ee;
        mem[237] = 10'h286;
        mem[238] = 10'h32a;
        mem[239] = 10'h067;
        mem[240] = 10'h2a2;
        mem[241] = 10'h1c3;
        mem[242] = 10'h126;
        mem[243] = 10'h0af;
        mem[244] = 10'h1e3;
        mem[245] = 10'h0ea;
        mem[246] = 10'h381;
        mem[247] = 10'h1f2;
        mem[248] = 10'h01a;
        mem[249] = 10'h1b2;
        mem[250] = 10'h215;
        mem[251] = 10'h36d;
        mem[252] = 10'h3ab;
        mem[253] = 10'h1cb;
        mem[254] = 10'h131;
        mem[255] = 10'h01c;
        mem[256] = 10'h0a9;
        mem[257] = 10'h369;
        mem[258] = 10'h096;
        mem[259] = 10'h2a1;
        mem[260] = 10'h070;
        mem[261] = 10'h196;
        mem[262] = 10'h0a8;
        mem[263] = 10'h3ed;
        mem[264] = 10'h071;
        mem[265] = 10'h2d7;
        mem[266] = 10'h0c7;
        mem[267] = 10'h28c;
        mem[268] = 10'h26e;
        mem[269] = 10'h0dd;
        mem[270] = 10'h010;
        mem[271] = 10'h140;
        mem[272] = 10'h159;
        mem[273] = 10'h19c;
        mem[274] = 10'h1a7;
        mem[275] = 10'h267;
        mem[276] = 10'h0ff;
        mem[277] = 10'h352;
        mem[278] = 10'h2ab;
        mem[279] = 10'h26d;
        mem[280] = 10'h362;
        mem[281] = 10'h24f;
        mem[282] = 10'h183;
        mem[283] = 10'h0cd;
        mem[284] = 10'h1c2;
        mem[285] = 10'h024;
        mem[286] = 10'h28b;
        mem[287] = 10'h206;
        mem[288] = 10'h1a9;
        mem[289] = 10'h0a2;
        mem[290] = 10'h016;
        mem[291] = 10'h34b;
        mem[292] = 10'h16f;
        mem[293] = 10'h2fd;
        mem[294] = 10'h0b6;
        mem[295] = 10'h2ff;
        mem[296] = 10'h242;
        mem[297] = 10'h0e6;
        mem[298] = 10'h2fe;
        mem[299] = 10'h1c6;
        mem[300] = 10'h1a4;
        mem[301] = 10'h17e;
        mem[302] = 10'h1a2;
        mem[303] = 10'h2d9;
        mem[304] = 10'h276;
        mem[305] = 10'h2fa;
        mem[306] = 10'h327;
        mem[307] = 10'h33b;
        mem[308] = 10'h243;
        mem[309] = 10'h3c8;
        mem[310] = 10'h05f;
        mem[311] = 10'h07d;
        mem[312] = 10'h07a;
        mem[313] = 10'h32f;
        mem[314] = 10'h009;
        mem[315] = 10'h3f3;
        mem[316] = 10'h09d;
        mem[317] = 10'h174;
        mem[318] = 10'h193;
        mem[319] = 10'h2bf;
        mem[320] = 10'h330;
        mem[321] = 10'h28d;
        mem[322] = 10'h3aa;
        mem[323] = 10'h068;
        mem[324] = 10'h333;
        mem[325] = 10'h1aa;
        mem[326] = 10'h356;
        mem[327] = 10'h2b3;
        mem[328] = 10'h3fe;
        mem[329] = 10'h007;
        mem[330] = 10'h2dd;
        mem[331] = 10'h2b0;
        mem[332] = 10'h3ae;
        mem[333] = 10'h12d;
        mem[334] = 10'h195;
        mem[335] = 10'h260;
        mem[336] = 10'h003;
        mem[337] = 10'h028;
        mem[338] = 10'h343;
        mem[339] = 10'h270;
        mem[340] = 10'h2d2;
        mem[341] = 10'h2cb;
        mem[342] = 10'h03b;
        mem[343] = 10'h218;
        mem[344] = 10'h16d;
        mem[345] = 10'h2eb;
        mem[346] = 10'h273;
        mem[347] = 10'h160;
        mem[348] = 10'h262;
        mem[349] = 10'h2be;
        mem[350] = 10'h143;
        mem[351] = 10'h0bd;
        mem[352] = 10'h27f;
        mem[353] = 10'h1c0;
        mem[354] = 10'h3e5;
        mem[355] = 10'h321;
        mem[356] = 10'h192;
        mem[357] = 10'h1c9;
        mem[358] = 10'h18d;
        mem[359] = 10'h142;
        mem[360] = 10'h0ae;
        mem[361] = 10'h237;
        mem[362] = 10'h037;
        mem[363] = 10'h0e3;
        mem[364] = 10'h3a3;
        mem[365] = 10'h389;
        mem[366] = 10'h2db;
        mem[367] = 10'h31d;
        mem[368] = 10'h07e;
        mem[369] = 10'h245;
        mem[370] = 10'h1c4;
        mem[371] = 10'h210;
        mem[372] = 10'h2a7;
        mem[373] = 10'h3e6;
        mem[374] = 10'h3f6;
        mem[375] = 10'h3de;
        mem[376] = 10'h344;
        mem[377] = 10'h325;
        mem[378] = 10'h399;
        mem[379] = 10'h034;
        mem[380] = 10'h172;
        mem[381] = 10'h251;
        mem[382] = 10'h2c6;
        mem[383] = 10'h130;
        mem[384] = 10'h15b;
        mem[385] = 10'h29e;
        mem[386] = 10'h305;
        mem[387] = 10'h3c5;
        mem[388] = 10'h27a;
        mem[389] = 10'h1a5;
        mem[390] = 10'h1fa;
        mem[391] = 10'h111;
        mem[392] = 10'h076;
        mem[393] = 10'h1c8;
        mem[394] = 10'h209;
        mem[395] = 10'h296;
        mem[396] = 10'h0e8;
        mem[397] = 10'h263;
        mem[398] = 10'h38a;
        mem[399] = 10'h050;
        mem[400] = 10'h004;
        mem[401] = 10'h31c;
        mem[402] = 10'h1f0;
        mem[403] = 10'h21f;
        mem[404] = 10'h048;
        mem[405] = 10'h379;
        mem[406] = 10'h141;
        mem[407] = 10'h015;
        mem[408] = 10'h39e;
        mem[409] = 10'h32d;
        mem[410] = 10'h323;
        mem[411] = 10'h25c;
        mem[412] = 10'h3f9;
        mem[413] = 10'h25f;
        mem[414] = 10'h315;
        mem[415] = 10'h34f;
        mem[416] = 10'h091;
        mem[417] = 10'h3c4;
        mem[418] = 10'h366;
        mem[419] = 10'h017;
        mem[420] = 10'h221;
        mem[421] = 10'h21d;
        mem[422] = 10'h17d;
        mem[423] = 10'h205;
        mem[424] = 10'h14b;
        mem[425] = 10'h0d0;
        mem[426] = 10'h3d9;
        mem[427] = 10'h291;
        mem[428] = 10'h04a;
        mem[429] = 10'h3c9;
        mem[430] = 10'h2e0;
        mem[431] = 10'h026;
        mem[432] = 10'h02a;
        mem[433] = 10'h3a0;
        mem[434] = 10'h00d;
        mem[435] = 10'h1f8;
        mem[436] = 10'h3cc;
        mem[437] = 10'h29c;
        mem[438] = 10'h08e;
        mem[439] = 10'h062;
        mem[440] = 10'h1ff;
        mem[441] = 10'h335;
        mem[442] = 10'h2b8;
        mem[443] = 10'h0cf;
        mem[444] = 10'h025;
        mem[445] = 10'h3e3;
        mem[446] = 10'h225;
        mem[447] = 10'h144;
        mem[448] = 10'h30b;
        mem[449] = 10'h2cd;
        mem[450] = 10'h22c;
        mem[451] = 10'h0c6;
        mem[452] = 10'h165;
        mem[453] = 10'h3bc;
        mem[454] = 10'h118;
        mem[455] = 10'h229;
        mem[456] = 10'h121;
        mem[457] = 10'h011;
        mem[458] = 10'h064;
        mem[459] = 10'h13c;
        mem[460] = 10'h16a;
        mem[461] = 10'h230;
        mem[462] = 10'h1e7;
        mem[463] = 10'h25d;
        mem[464] = 10'h329;
        mem[465] = 10'h00c;
        mem[466] = 10'h02f;
        mem[467] = 10'h17b;
        mem[468] = 10'h26f;
        mem[469] = 10'h188;
        mem[470] = 10'h042;
        mem[471] = 10'h164;
        mem[472] = 10'h0d2;
        mem[473] = 10'h30a;
        mem[474] = 10'h109;
        mem[475] = 10'h306;
        mem[476] = 10'h018;
        mem[477] = 10'h1e9;
        mem[478] = 10'h059;
        mem[479] = 10'h1f1;
        mem[480] = 10'h0ba;
        mem[481] = 10'h281;
        mem[482] = 10'h058;
        mem[483] = 10'h081;
        mem[484] = 10'h2d1;
        mem[485] = 10'h057;
        mem[486] = 10'h0e2;
        mem[487] = 10'h2d0;
        mem[488] = 10'h1cd;
        mem[489] = 10'h375;
        mem[490] = 10'h254;
        mem[491] = 10'h2cc;
        mem[492] = 10'h178;
        mem[493] = 10'h363;
        mem[494] = 10'h1a6;
        mem[495] = 10'h32b;
        mem[496] = 10'h226;
        mem[497] = 10'h204;
        mem[498] = 10'h359;
        mem[499] = 10'h22d;
        mem[500] = 10'h3b9;
        mem[501] = 10'h0b9;
        mem[502] = 10'h044;
        mem[503] = 10'h1fe;
        mem[504] = 10'h23c;
        mem[505] = 10'h3b8;
        mem[506] = 10'h1c5;
        mem[507] = 10'h34d;
        mem[508] = 10'h1ac;
        mem[509] = 10'h355;
        mem[510] = 10'h1e1;
        mem[511] = 10'h006;
        mem[512] = 10'h1b0;
        mem[513] = 10'h280;
        mem[514] = 10'h1ed;
        mem[515] = 10'h098;
        mem[516] = 10'h284;
        mem[517] = 10'h05d;
        mem[518] = 10'h030;
        mem[519] = 10'h23e;
        mem[520] = 10'h092;
        mem[521] = 10'h134;
        mem[522] = 10'h1fb;
        mem[523] = 10'h2aa;
        mem[524] = 10'h043;
        mem[525] = 10'h1b7;
        mem[526] = 10'h2e4;
        mem[527] = 10'h021;
        mem[528] = 10'h388;
        mem[529] = 10'h3dd;
        mem[530] = 10'h10c;
        mem[531] = 10'h309;
        mem[532] = 10'h145;
        mem[533] = 10'h35c;
        mem[534] = 10'h1cc;
        mem[535] = 10'h00f;
        mem[536] = 10'h18c;
        mem[537] = 10'h056;
        mem[538] = 10'h146;
        mem[539] = 10'h2b4;
        mem[540] = 10'h171;
        mem[541] = 10'h3f0;
        mem[542] = 10'h14f;
        mem[543] = 10'h027;
        mem[544] = 10'h1ce;
        mem[545] = 10'h06d;
        mem[546] = 10'h38c;
        mem[547] = 10'h1c7;
        mem[548] = 10'h378;
        mem[549] = 10'h36c;
        mem[550] = 10'h0e5;
        mem[551] = 10'h3f2;
        mem[552] = 10'h0b2;
        mem[553] = 10'h211;
        mem[554] = 10'h19f;
        mem[555] = 10'h308;
        mem[556] = 10'h14d;
        mem[557] = 10'h069;
        mem[558] = 10'h3b7;
        mem[559] = 10'h256;
        mem[560] = 10'h2a8;
        mem[561] = 10'h353;
        mem[562] = 10'h116;
        mem[563] = 10'h3ef;
        mem[564] = 10'h082;
        mem[565] = 10'h3c2;
        mem[566] = 10'h2bb;
        mem[567] = 10'h2df;
        mem[568] = 10'h0a4;
        mem[569] = 10'h167;
        mem[570] = 10'h392;
        mem[571] = 10'h29a;
        mem[572] = 10'h0c4;
        mem[573] = 10'h3ea;
        mem[574] = 10'h0b4;
        mem[575] = 10'h20c;
        mem[576] = 10'h2ad;
        mem[577] = 10'h3fb;
        mem[578] = 10'h180;
        mem[579] = 10'h19e;
        mem[580] = 10'h087;
        mem[581] = 10'h37d;
        mem[582] = 10'h36b;
        mem[583] = 10'h14c;
        mem[584] = 10'h1da;
        mem[585] = 10'h0d9;
        mem[586] = 10'h0e1;
        mem[587] = 10'h0bf;
        mem[588] = 10'h2af;
        mem[589] = 10'h1d4;
        mem[590] = 10'h334;
        mem[591] = 10'h094;
        mem[592] = 10'h114;
        mem[593] = 10'h3ad;
        mem[594] = 10'h2d4;
        mem[595] = 10'h3ca;
        mem[596] = 10'h03a;
        mem[597] = 10'h2b1;
        mem[598] = 10'h0b8;
        mem[599] = 10'h1dc;
        mem[600] = 10'h2f5;
        mem[601] = 10'h214;
        mem[602] = 10'h25b;
        mem[603] = 10'h2a0;
        mem[604] = 10'h35d;
        mem[605] = 10'h2c0;
        mem[606] = 10'h3c0;
        mem[607] = 10'h33e;
        mem[608] = 10'h27c;
        mem[609] = 10'h37e;
        mem[610] = 10'h0cb;
        mem[611] = 10'h0d1;
        mem[612] = 10'h247;
        mem[613] = 10'h005;
        mem[614] = 10'h1f3;
        mem[615] = 10'h36e;
        mem[616] = 10'h224;
        mem[617] = 10'h0de;
        mem[618] = 10'h3f7;
        mem[619] = 10'h122;
        mem[620] = 10'h13d;
        mem[621] = 10'h37b;
        mem[622] = 10'h17f;
        mem[623] = 10'h396;
        mem[624] = 10'h32c;
        mem[625] = 10'h184;
        mem[626] = 10'h1e8;
        mem[627] = 10'h1b3;
        mem[628] = 10'h35b;
        mem[629] = 10'h259;
        mem[630] = 10'h269;
        mem[631] = 10'h182;
        mem[632] = 10'h1df;
        mem[633] = 10'h18a;
        mem[634] = 10'h2f3;
        mem[635] = 10'h33d;
        mem[636] = 10'h301;
        mem[637] = 10'h033;
        mem[638] = 10'h21a;
        mem[639] = 10'h19a;
        mem[640] = 10'h199;
        mem[641] = 10'h0c9;
        mem[642] = 10'h223;
        mem[643] = 10'h039;
        mem[644] = 10'h0fd;
        mem[645] = 10'h30d;
        mem[646] = 10'h24d;
        mem[647] = 10'h055;
        mem[648] = 10'h150;
        mem[649] = 10'h385;
        mem[650] = 10'h1ea;
        mem[651] = 10'h2c7;
        mem[652] = 10'h04f;
        mem[653] = 10'h266;
        mem[654] = 10'h1d5;
        mem[655] = 10'h1d0;
        mem[656] = 10'h22f;
        mem[657] = 10'h089;
        mem[658] = 10'h102;
        mem[659] = 10'h105;
        mem[660] = 10'h23d;
        mem[661] = 10'h30e;
        mem[662] = 10'h0f3;
        mem[663] = 10'h15e;
        mem[664] = 10'h038;
        mem[665] = 10'h124;
        mem[666] = 10'h132;
        mem[667] = 10'h019;
        mem[668] = 10'h3c6;
        mem[669] = 10'h324;
        mem[670] = 10'h3a2;
        mem[671] = 10'h162;
        mem[672] = 10'h2bd;
        mem[673] = 10'h1eb;
        mem[674] = 10'h138;
        mem[675] = 10'h08d;
        mem[676] = 10'h22b;
        mem[677] = 10'h2bc;
        mem[678] = 10'h176;
        mem[679] = 10'h041;
        mem[680] = 10'h2c1;
        mem[681] = 10'h3bf;
        mem[682] = 10'h24c;
        mem[683] = 10'h3d7;
        mem[684] = 10'h0b1;
        mem[685] = 10'h24b;
        mem[686] = 10'h3fd;
        mem[687] = 10'h0f4;
        mem[688] = 10'h052;
        mem[689] = 10'h100;
        mem[690] = 10'h2ea;
        mem[691] = 10'h0dc;
        mem[692] = 10'h2ed;
        mem[693] = 10'h2b2;
        mem[694] = 10'h1f5;
        mem[695] = 10'h257;
        mem[696] = 10'h2f2;
        mem[697] = 10'h21c;
        mem[698] = 10'h2f6;
        mem[699] = 10'h0fc;
        mem[700] = 10'h374;
        mem[701] = 10'h289;
        mem[702] = 10'h086;
        mem[703] = 10'h0e7;
        mem[704] = 10'h233;
        mem[705] = 10'h3e7;
        mem[706] = 10'h1b4;
        mem[707] = 10'h1ae;
        mem[708] = 10'h07f;
        mem[709] = 10'h2e2;
        mem[710] = 10'h19d;
        mem[711] = 10'h365;
        mem[712] = 10'h371;
        mem[713] = 10'h342;
        mem[714] = 10'h1d2;
        mem[715] = 10'h11b;
        mem[716] = 10'h3f8;
        mem[717] = 10'h1f7;
        mem[718] = 10'h38e;
        mem[719] = 10'h2a6;
        mem[720] = 10'h17a;
        mem[721] = 10'h2c4;
        mem[722] = 10'h20e;
        mem[723] = 10'h1bd;
        mem[724] = 10'h312;
        mem[725] = 10'h09c;
        mem[726] = 10'h000;
        mem[727] = 10'h240;
        mem[728] = 10'h2de;
        mem[729] = 10'h26c;
        mem[730] = 10'h10a;
        mem[731] = 10'h11d;
        mem[732] = 10'h231;
        mem[733] = 10'h382;
        mem[734] = 10'h0aa;
        mem[735] = 10'h19b;
        mem[736] = 10'h370;
        mem[737] = 10'h398;
        mem[738] = 10'h31b;
        mem[739] = 10'h2e7;
        mem[740] = 10'h300;
        mem[741] = 10'h3b5;
        mem[742] = 10'h014;
        mem[743] = 10'h093;
        mem[744] = 10'h103;
        mem[745] = 10'h319;
        mem[746] = 10'h1a3;
        mem[747] = 10'h2b9;
        mem[748] = 10'h173;
        mem[749] = 10'h3cd;
        mem[750] = 10'h1b9;
        mem[751] = 10'h03f;
        mem[752] = 10'h0d5;
        mem[753] = 10'h09b;
        mem[754] = 10'h3ba;
        mem[755] = 10'h084;
        mem[756] = 10'h127;
        mem[757] = 10'h0b7;
        mem[758] = 10'h339;
        mem[759] = 10'h1e0;
        mem[760] = 10'h03c;
        mem[761] = 10'h3a5;
        mem[762] = 10'h077;
        mem[763] = 10'h3e1;
        mem[764] = 10'h1c1;
        mem[765] = 10'h3e0;
        mem[766] = 10'h002;
        mem[767] = 10'h18f;
        mem[768] = 10'h106;
        mem[769] = 10'h0c2;
        mem[770] = 10'h1fd;
        mem[771] = 10'h179;
        mem[772] = 10'h0d8;
        mem[773] = 10'h3bb;
        mem[774] = 10'h2a5;
        mem[775] = 10'h39d;
        mem[776] = 10'h258;
        mem[777] = 10'h28f;
        mem[778] = 10'h328;
        mem[779] = 10'h0ec;
        mem[780] = 10'h3d1;
        mem[781] = 10'h168;
        mem[782] = 10'h3d8;
        mem[783] = 10'h045;
        mem[784] = 10'h26b;
        mem[785] = 10'h0f2;
        mem[786] = 10'h123;
        mem[787] = 10'h060;
        mem[788] = 10'h0b5;
        mem[789] = 10'h39a;
        mem[790] = 10'h27e;
        mem[791] = 10'h307;
        mem[792] = 10'h190;
        mem[793] = 10'h2e9;
        mem[794] = 10'h239;
        mem[795] = 10'h09f;
        mem[796] = 10'h2a4;
        mem[797] = 10'h0bb;
        mem[798] = 10'h347;
        mem[799] = 10'h377;
        mem[800] = 10'h373;
        mem[801] = 10'h0e9;
        mem[802] = 10'h198;
        mem[803] = 10'h3b6;
        mem[804] = 10'h3e8;
        mem[805] = 10'h155;
        mem[806] = 10'h350;
        mem[807] = 10'h1b1;
        mem[808] = 10'h3d3;
        mem[809] = 10'h331;
        mem[810] = 10'h387;
        mem[811] = 10'h189;
        mem[812] = 10'h3ec;
        mem[813] = 10'h21b;
        mem[814] = 10'h351;
        mem[815] = 10'h1af;
        mem[816] = 10'h3c3;
        mem[817] = 10'h049;
        mem[818] = 10'h393;
        mem[819] = 10'h2d8;
        mem[820] = 10'h0f1;
        mem[821] = 10'h292;
        mem[822] = 10'h0d6;
        mem[823] = 10'h35a;
        mem[824] = 10'h332;
        mem[825] = 10'h235;
        mem[826] = 10'h22e;
        mem[827] = 10'h28a;
        mem[828] = 10'h0d7;
        mem[829] = 10'h386;
        mem[830] = 10'h02d;
        mem[831] = 10'h00b;
        mem[832] = 10'h097;
        mem[833] = 10'h310;
        mem[834] = 10'h29d;
        mem[835] = 10'h3f1;
        mem[836] = 10'h09a;
        mem[837] = 10'h2f8;
        mem[838] = 10'h31e;
        mem[839] = 10'h349;
        mem[840] = 10'h3d6;
        mem[841] = 10'h391;
        mem[842] = 10'h0c0;
        mem[843] = 10'h228;
        mem[844] = 10'h1d7;
        mem[845] = 10'h012;
        mem[846] = 10'h07c;
        mem[847] = 10'h1f9;
        mem[848] = 10'h299;
        mem[849] = 10'h354;
        mem[850] = 10'h271;
        mem[851] = 10'h083;
        mem[852] = 10'h11c;
        mem[853] = 10'h0d4;
        mem[854] = 10'h23f;
        mem[855] = 10'h0f8;
        mem[856] = 10'h151;
        mem[857] = 10'h108;
        mem[858] = 10'h203;
        mem[859] = 10'h181;
        mem[860] = 10'h3fc;
        mem[861] = 10'h217;
        mem[862] = 10'h3e9;
        mem[863] = 10'h163;
        mem[864] = 10'h107;
        mem[865] = 10'h12b;
        mem[866] = 10'h232;
        mem[867] = 10'h2f0;
        mem[868] = 10'h166;
        mem[869] = 10'h394;
        mem[870] = 10'h0bc;
        mem[871] = 10'h38b;
        mem[872] = 10'h288;
        mem[873] = 10'h287;
        mem[874] = 10'h3a4;
        mem[875] = 10'h175;
        mem[876] = 10'h15c;
        mem[877] = 10'h0cc;
        mem[878] = 10'h136;
        mem[879] = 10'h3cb;
        mem[880] = 10'h208;
        mem[881] = 10'h338;
        mem[882] = 10'h0fa;
        mem[883] = 10'h10d;
        mem[884] = 10'h16c;
        mem[885] = 10'h2d6;
        mem[886] = 10'h0da;
        mem[887] = 10'h1a8;
        mem[888] = 10'h361;
        mem[889] = 10'h0ac;
        mem[890] = 10'h187;
        mem[891] = 10'h249;
        mem[892] = 10'h022;
        mem[893] = 10'h1d6;
        mem[894] = 10'h08f;
        mem[895] = 10'h065;
        mem[896] = 10'h156;
        mem[897] = 10'h0f7;
        mem[898] = 10'h3a6;
        mem[899] = 10'h3b1;
        mem[900] = 10'h3a1;
        mem[901] = 10'h29f;
        mem[902] = 10'h1ec;
        mem[903] = 10'h0db;
        mem[904] = 10'h061;
        mem[905] = 10'h0c5;
        mem[906] = 10'h0be;
        mem[907] = 10'h133;
        mem[908] = 10'h13a;
        mem[909] = 10'h20d;
        mem[910] = 10'h013;
        mem[911] = 10'h2e1;
        mem[912] = 10'h1f4;
        mem[913] = 10'h318;
        mem[914] = 10'h1de;
        mem[915] = 10'h12f;
        mem[916] = 10'h30c;
        mem[917] = 10'h2e6;
        mem[918] = 10'h201;
        mem[919] = 10'h397;
        mem[920] = 10'h0f9;
        mem[921] = 10'h384;
        mem[922] = 10'h115;
        mem[923] = 10'h2a3;
        mem[924] = 10'h2e3;
        mem[925] = 10'h336;
        mem[926] = 10'h364;
        mem[927] = 10'h295;
        mem[928] = 10'h0a1;
        mem[929] = 10'h11a;
        mem[930] = 10'h169;
        mem[931] = 10'h047;
        mem[932] = 10'h0b0;
        mem[933] = 10'h2c9;
        mem[934] = 10'h248;
        mem[935] = 10'h1cf;
        mem[936] = 10'h05a;
        mem[937] = 10'h37f;
        mem[938] = 10'h0fe;
        mem[939] = 10'h238;
        mem[940] = 10'h2c8;
        mem[941] = 10'h03e;
        mem[942] = 10'h3dc;
        mem[943] = 10'h16b;
        mem[944] = 10'h341;
        mem[945] = 10'h0f5;
        mem[946] = 10'h16e;
        mem[947] = 10'h2a9;
        mem[948] = 10'h080;
        mem[949] = 10'h1e5;
        mem[950] = 10'h297;
        mem[951] = 10'h1ba;
        mem[952] = 10'h154;
        mem[953] = 10'h253;
        mem[954] = 10'h18b;
        mem[955] = 10'h119;
        mem[956] = 10'h34e;
        mem[957] = 10'h008;
        mem[958] = 10'h158;
        mem[959] = 10'h261;
        mem[960] = 10'h0ce;
        mem[961] = 10'h148;
        mem[962] = 10'h33c;
        mem[963] = 10'h2f4;
        mem[964] = 10'h05e;
        mem[965] = 10'h30f;
        mem[966] = 10'h24a;
        mem[967] = 10'h255;
        mem[968] = 10'h3ce;
        mem[969] = 10'h234;
        mem[970] = 10'h2e8;
        mem[971] = 10'h0ab;
        mem[972] = 10'h3b3;
        mem[973] = 10'h0a5;
        mem[974] = 10'h02c;
        mem[975] = 10'h304;
        mem[976] = 10'h294;
        mem[977] = 10'h01d;
        mem[978] = 10'h348;
        mem[979] = 10'h0a7;
        mem[980] = 10'h15f;
        mem[981] = 10'h275;
        mem[982] = 10'h36f;
        mem[983] = 10'h1fc;
        mem[984] = 10'h1ca;
        mem[985] = 10'h3c1;
        mem[986] = 10'h10e;
        mem[987] = 10'h1e2;
        mem[988] = 10'h01b;
        mem[989] = 10'h2b5;
        mem[990] = 10'h066;
        mem[991] = 10'h360;
        mem[992] = 10'h265;
        mem[993] = 10'h268;
        mem[994] = 10'h33f;
        mem[995] = 10'h11f;
        mem[996] = 10'h326;
        mem[997] = 10'h1d1;
        mem[998] = 10'h08b;
        mem[999] = 10'h345;
        mem[1000] = 10'h2e5;
        mem[1001] = 10'h340;
        mem[1002] = 10'h1bc;
        mem[1003] = 10'h3f4;
        mem[1004] = 10'h3d5;
        mem[1005] = 10'h088;
        mem[1006] = 10'h18e;
        mem[1007] = 10'h279;
        mem[1008] = 10'h3bd;
        mem[1009] = 10'h2ba;
        mem[1010] = 10'h283;
        mem[1011] = 10'h06a;
        mem[1012] = 10'h2ae;
        mem[1013] = 10'h202;
        mem[1014] = 10'h02e;
        mem[1015] = 10'h2ca;
        mem[1016] = 10'h117;
        mem[1017] = 10'h35f;
        mem[1018] = 10'h322;
        mem[1019] = 10'h2c2;
        mem[1020] = 10'h14a;
        mem[1021] = 10'h320;
        mem[1022] = 10'h395;
        mem[1023] = 10'h2c3;
    end
endmodule

module encrypt_4sbox_large5(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h2d3;
        mem[1] = 10'h325;
        mem[2] = 10'h1f0;
        mem[3] = 10'h007;
        mem[4] = 10'h396;
        mem[5] = 10'h04f;
        mem[6] = 10'h35b;
        mem[7] = 10'h24e;
        mem[8] = 10'h21d;
        mem[9] = 10'h287;
        mem[10] = 10'h178;
        mem[11] = 10'h18d;
        mem[12] = 10'h32f;
        mem[13] = 10'h16e;
        mem[14] = 10'h0f8;
        mem[15] = 10'h3ce;
        mem[16] = 10'h3ab;
        mem[17] = 10'h31a;
        mem[18] = 10'h24c;
        mem[19] = 10'h2c9;
        mem[20] = 10'h343;
        mem[21] = 10'h179;
        mem[22] = 10'h24a;
        mem[23] = 10'h1a0;
        mem[24] = 10'h223;
        mem[25] = 10'h26d;
        mem[26] = 10'h208;
        mem[27] = 10'h308;
        mem[28] = 10'h260;
        mem[29] = 10'h242;
        mem[30] = 10'h267;
        mem[31] = 10'h317;
        mem[32] = 10'h10b;
        mem[33] = 10'h246;
        mem[34] = 10'h385;
        mem[35] = 10'h168;
        mem[36] = 10'h19b;
        mem[37] = 10'h189;
        mem[38] = 10'h03a;
        mem[39] = 10'h19d;
        mem[40] = 10'h2aa;
        mem[41] = 10'h1b4;
        mem[42] = 10'h39f;
        mem[43] = 10'h1a5;
        mem[44] = 10'h2eb;
        mem[45] = 10'h139;
        mem[46] = 10'h0af;
        mem[47] = 10'h09f;
        mem[48] = 10'h0c3;
        mem[49] = 10'h3cc;
        mem[50] = 10'h371;
        mem[51] = 10'h0f0;
        mem[52] = 10'h01c;
        mem[53] = 10'h39e;
        mem[54] = 10'h0f9;
        mem[55] = 10'h33d;
        mem[56] = 10'h23b;
        mem[57] = 10'h11c;
        mem[58] = 10'h0f7;
        mem[59] = 10'h324;
        mem[60] = 10'h227;
        mem[61] = 10'h355;
        mem[62] = 10'h2a4;
        mem[63] = 10'h3f4;
        mem[64] = 10'h101;
        mem[65] = 10'h0fe;
        mem[66] = 10'h2c7;
        mem[67] = 10'h330;
        mem[68] = 10'h12b;
        mem[69] = 10'h205;
        mem[70] = 10'h063;
        mem[71] = 10'h273;
        mem[72] = 10'h2bb;
        mem[73] = 10'h38c;
        mem[74] = 10'h1fa;
        mem[75] = 10'h07d;
        mem[76] = 10'h100;
        mem[77] = 10'h251;
        mem[78] = 10'h18b;
        mem[79] = 10'h22b;
        mem[80] = 10'h01b;
        mem[81] = 10'h049;
        mem[82] = 10'h3d6;
        mem[83] = 10'h1e0;
        mem[84] = 10'h214;
        mem[85] = 10'h284;
        mem[86] = 10'h156;
        mem[87] = 10'h30d;
        mem[88] = 10'h15a;
        mem[89] = 10'h05d;
        mem[90] = 10'h376;
        mem[91] = 10'h22f;
        mem[92] = 10'h390;
        mem[93] = 10'h00e;
        mem[94] = 10'h3a0;
        mem[95] = 10'h2b5;
        mem[96] = 10'h040;
        mem[97] = 10'h027;
        mem[98] = 10'h2b4;
        mem[99] = 10'h1f7;
        mem[100] = 10'h1f4;
        mem[101] = 10'h00d;
        mem[102] = 10'h3fa;
        mem[103] = 10'h00f;
        mem[104] = 10'h2a0;
        mem[105] = 10'h259;
        mem[106] = 10'h2ac;
        mem[107] = 10'h3d2;
        mem[108] = 10'h191;
        mem[109] = 10'h33c;
        mem[110] = 10'h2e4;
        mem[111] = 10'h0d1;
        mem[112] = 10'h3ae;
        mem[113] = 10'h337;
        mem[114] = 10'h07e;
        mem[115] = 10'h3ba;
        mem[116] = 10'h0a1;
        mem[117] = 10'h04d;
        mem[118] = 10'h3fe;
        mem[119] = 10'h31e;
        mem[120] = 10'h30c;
        mem[121] = 10'h076;
        mem[122] = 10'h297;
        mem[123] = 10'h008;
        mem[124] = 10'h3a6;
        mem[125] = 10'h084;
        mem[126] = 10'h2b3;
        mem[127] = 10'h2bf;
        mem[128] = 10'h217;
        mem[129] = 10'h204;
        mem[130] = 10'h2fb;
        mem[131] = 10'h1ff;
        mem[132] = 10'h269;
        mem[133] = 10'h20e;
        mem[134] = 10'h1af;
        mem[135] = 10'h25c;
        mem[136] = 10'h1f8;
        mem[137] = 10'h186;
        mem[138] = 10'h0ab;
        mem[139] = 10'h0df;
        mem[140] = 10'h13f;
        mem[141] = 10'h1e1;
        mem[142] = 10'h046;
        mem[143] = 10'h3ec;
        mem[144] = 10'h202;
        mem[145] = 10'h1c2;
        mem[146] = 10'h1e2;
        mem[147] = 10'h3c0;
        mem[148] = 10'h16a;
        mem[149] = 10'h27b;
        mem[150] = 10'h021;
        mem[151] = 10'h314;
        mem[152] = 10'h228;
        mem[153] = 10'h1e7;
        mem[154] = 10'h3db;
        mem[155] = 10'h194;
        mem[156] = 10'h2a5;
        mem[157] = 10'h03d;
        mem[158] = 10'h200;
        mem[159] = 10'h0fc;
        mem[160] = 10'h203;
        mem[161] = 10'h2f2;
        mem[162] = 10'h08d;
        mem[163] = 10'h257;
        mem[164] = 10'h264;
        mem[165] = 10'h306;
        mem[166] = 10'h3bc;
        mem[167] = 10'h10c;
        mem[168] = 10'h249;
        mem[169] = 10'h001;
        mem[170] = 10'h2cd;
        mem[171] = 10'h350;
        mem[172] = 10'h1d3;
        mem[173] = 10'h0b3;
        mem[174] = 10'h3cf;
        mem[175] = 10'h258;
        mem[176] = 10'h231;
        mem[177] = 10'h11d;
        mem[178] = 10'h239;
        mem[179] = 10'h211;
        mem[180] = 10'h03e;
        mem[181] = 10'h309;
        mem[182] = 10'h0d3;
        mem[183] = 10'h3ef;
        mem[184] = 10'h340;
        mem[185] = 10'h393;
        mem[186] = 10'h20f;
        mem[187] = 10'h0bc;
        mem[188] = 10'h17f;
        mem[189] = 10'h2af;
        mem[190] = 10'h37c;
        mem[191] = 10'h379;
        mem[192] = 10'h1eb;
        mem[193] = 10'h232;
        mem[194] = 10'h094;
        mem[195] = 10'h3d9;
        mem[196] = 10'h1ba;
        mem[197] = 10'h25a;
        mem[198] = 10'h1f5;
        mem[199] = 10'h2ae;
        mem[200] = 10'h1d0;
        mem[201] = 10'h336;
        mem[202] = 10'h187;
        mem[203] = 10'h0c8;
        mem[204] = 10'h079;
        mem[205] = 10'h256;
        mem[206] = 10'h096;
        mem[207] = 10'h1a6;
        mem[208] = 10'h068;
        mem[209] = 10'h04e;
        mem[210] = 10'h1f9;
        mem[211] = 10'h29c;
        mem[212] = 10'h17b;
        mem[213] = 10'h134;
        mem[214] = 10'h11f;
        mem[215] = 10'h059;
        mem[216] = 10'h347;
        mem[217] = 10'h1d6;
        mem[218] = 10'h044;
        mem[219] = 10'h0e5;
        mem[220] = 10'h0bf;
        mem[221] = 10'h07b;
        mem[222] = 10'h0e4;
        mem[223] = 10'h031;
        mem[224] = 10'h2dd;
        mem[225] = 10'h0e0;
        mem[226] = 10'h3ca;
        mem[227] = 10'h3a2;
        mem[228] = 10'h0c6;
        mem[229] = 10'h345;
        mem[230] = 10'h23f;
        mem[231] = 10'h31b;
        mem[232] = 10'h3a9;
        mem[233] = 10'h279;
        mem[234] = 10'h233;
        mem[235] = 10'h02c;
        mem[236] = 10'h277;
        mem[237] = 10'h14f;
        mem[238] = 10'h1fe;
        mem[239] = 10'h2a3;
        mem[240] = 10'h2f5;
        mem[241] = 10'h3ed;
        mem[242] = 10'h092;
        mem[243] = 10'h352;
        mem[244] = 10'h2b2;
        mem[245] = 10'h1ee;
        mem[246] = 10'h365;
        mem[247] = 10'h20d;
        mem[248] = 10'h015;
        mem[249] = 10'h263;
        mem[250] = 10'h032;
        mem[251] = 10'h266;
        mem[252] = 10'h1c9;
        mem[253] = 10'h36e;
        mem[254] = 10'h2de;
        mem[255] = 10'h1cf;
        mem[256] = 10'h210;
        mem[257] = 10'h3aa;
        mem[258] = 10'h23d;
        mem[259] = 10'h3b1;
        mem[260] = 10'h234;
        mem[261] = 10'h08e;
        mem[262] = 10'h1c1;
        mem[263] = 10'h143;
        mem[264] = 10'h3a4;
        mem[265] = 10'h3cd;
        mem[266] = 10'h2c1;
        mem[267] = 10'h017;
        mem[268] = 10'h302;
        mem[269] = 10'h3b8;
        mem[270] = 10'h34d;
        mem[271] = 10'h0ee;
        mem[272] = 10'h0ed;
        mem[273] = 10'h1ac;
        mem[274] = 10'h1c7;
        mem[275] = 10'h26a;
        mem[276] = 10'h383;
        mem[277] = 10'h169;
        mem[278] = 10'h262;
        mem[279] = 10'h3a3;
        mem[280] = 10'h299;
        mem[281] = 10'h368;
        mem[282] = 10'h061;
        mem[283] = 10'h11b;
        mem[284] = 10'h0a3;
        mem[285] = 10'h1d9;
        mem[286] = 10'h37f;
        mem[287] = 10'h0f6;
        mem[288] = 10'h248;
        mem[289] = 10'h2c0;
        mem[290] = 10'h1db;
        mem[291] = 10'h066;
        mem[292] = 10'h3c6;
        mem[293] = 10'h114;
        mem[294] = 10'h2ff;
        mem[295] = 10'h135;
        mem[296] = 10'h384;
        mem[297] = 10'h3af;
        mem[298] = 10'h133;
        mem[299] = 10'h38d;
        mem[300] = 10'h216;
        mem[301] = 10'h08c;
        mem[302] = 10'h2e3;
        mem[303] = 10'h36a;
        mem[304] = 10'h1e3;
        mem[305] = 10'h0c4;
        mem[306] = 10'h387;
        mem[307] = 10'h126;
        mem[308] = 10'h019;
        mem[309] = 10'h3b9;
        mem[310] = 10'h33b;
        mem[311] = 10'h075;
        mem[312] = 10'h138;
        mem[313] = 10'h270;
        mem[314] = 10'h3f1;
        mem[315] = 10'h13c;
        mem[316] = 10'h0ba;
        mem[317] = 10'h1e5;
        mem[318] = 10'h1ab;
        mem[319] = 10'h334;
        mem[320] = 10'h01e;
        mem[321] = 10'h1aa;
        mem[322] = 10'h0ae;
        mem[323] = 10'h243;
        mem[324] = 10'h35d;
        mem[325] = 10'h2d4;
        mem[326] = 10'h386;
        mem[327] = 10'h174;
        mem[328] = 10'h300;
        mem[329] = 10'h3e2;
        mem[330] = 10'h2c5;
        mem[331] = 10'h17d;
        mem[332] = 10'h1b7;
        mem[333] = 10'h1b1;
        mem[334] = 10'h160;
        mem[335] = 10'h394;
        mem[336] = 10'h2ee;
        mem[337] = 10'h2d6;
        mem[338] = 10'h07a;
        mem[339] = 10'h3e4;
        mem[340] = 10'h24f;
        mem[341] = 10'h1d1;
        mem[342] = 10'h060;
        mem[343] = 10'h0cc;
        mem[344] = 10'h261;
        mem[345] = 10'h28c;
        mem[346] = 10'h006;
        mem[347] = 10'h275;
        mem[348] = 10'h026;
        mem[349] = 10'h235;
        mem[350] = 10'h247;
        mem[351] = 10'h131;
        mem[352] = 10'h0a7;
        mem[353] = 10'h0cf;
        mem[354] = 10'h315;
        mem[355] = 10'h377;
        mem[356] = 10'h3e3;
        mem[357] = 10'h2fe;
        mem[358] = 10'h2b0;
        mem[359] = 10'h0cb;
        mem[360] = 10'h35a;
        mem[361] = 10'h167;
        mem[362] = 10'h10e;
        mem[363] = 10'h130;
        mem[364] = 10'h1ae;
        mem[365] = 10'h323;
        mem[366] = 10'h33a;
        mem[367] = 10'h0d7;
        mem[368] = 10'h184;
        mem[369] = 10'h225;
        mem[370] = 10'h29b;
        mem[371] = 10'h000;
        mem[372] = 10'h378;
        mem[373] = 10'h2ec;
        mem[374] = 10'h318;
        mem[375] = 10'h0e1;
        mem[376] = 10'h240;
        mem[377] = 10'h3c4;
        mem[378] = 10'h1f6;
        mem[379] = 10'h190;
        mem[380] = 10'h052;
        mem[381] = 10'h14b;
        mem[382] = 10'h0ac;
        mem[383] = 10'h3d1;
        mem[384] = 10'h0cd;
        mem[385] = 10'h2e8;
        mem[386] = 10'h17a;
        mem[387] = 10'h0d6;
        mem[388] = 10'h392;
        mem[389] = 10'h109;
        mem[390] = 10'h0b5;
        mem[391] = 10'h0a2;
        mem[392] = 10'h3c7;
        mem[393] = 10'h31f;
        mem[394] = 10'h1a7;
        mem[395] = 10'h20c;
        mem[396] = 10'h3b6;
        mem[397] = 10'h2ad;
        mem[398] = 10'h09a;
        mem[399] = 10'h082;
        mem[400] = 10'h3a1;
        mem[401] = 10'h3b7;
        mem[402] = 10'h36f;
        mem[403] = 10'h39c;
        mem[404] = 10'h2bc;
        mem[405] = 10'h177;
        mem[406] = 10'h2a8;
        mem[407] = 10'h3e0;
        mem[408] = 10'h37d;
        mem[409] = 10'h3fd;
        mem[410] = 10'h2e5;
        mem[411] = 10'h2a9;
        mem[412] = 10'h0f4;
        mem[413] = 10'h2e1;
        mem[414] = 10'h0e8;
        mem[415] = 10'h375;
        mem[416] = 10'h074;
        mem[417] = 10'h07c;
        mem[418] = 10'h30b;
        mem[419] = 10'h2f3;
        mem[420] = 10'h158;
        mem[421] = 10'h2c6;
        mem[422] = 10'h0c0;
        mem[423] = 10'h0b8;
        mem[424] = 10'h064;
        mem[425] = 10'h332;
        mem[426] = 10'h2e2;
        mem[427] = 10'h25e;
        mem[428] = 10'h0b1;
        mem[429] = 10'h182;
        mem[430] = 10'h0c5;
        mem[431] = 10'h3f5;
        mem[432] = 10'h1ef;
        mem[433] = 10'h02d;
        mem[434] = 10'h1a8;
        mem[435] = 10'h1c0;
        mem[436] = 10'h2b6;
        mem[437] = 10'h03b;
        mem[438] = 10'h1b2;
        mem[439] = 10'h21e;
        mem[440] = 10'h32e;
        mem[441] = 10'h1c3;
        mem[442] = 10'h2f1;
        mem[443] = 10'h29e;
        mem[444] = 10'h19f;
        mem[445] = 10'h33f;
        mem[446] = 10'h198;
        mem[447] = 10'h3be;
        mem[448] = 10'h1ed;
        mem[449] = 10'h12f;
        mem[450] = 10'h011;
        mem[451] = 10'h0dc;
        mem[452] = 10'h15b;
        mem[453] = 10'h3bb;
        mem[454] = 10'h305;
        mem[455] = 10'h2bd;
        mem[456] = 10'h1bc;
        mem[457] = 10'h27a;
        mem[458] = 10'h095;
        mem[459] = 10'h06f;
        mem[460] = 10'h3cb;
        mem[461] = 10'h3c9;
        mem[462] = 10'h022;
        mem[463] = 10'h1ca;
        mem[464] = 10'h09c;
        mem[465] = 10'h3ea;
        mem[466] = 10'h057;
        mem[467] = 10'h06d;
        mem[468] = 10'h311;
        mem[469] = 10'h3f7;
        mem[470] = 10'h2ab;
        mem[471] = 10'h151;
        mem[472] = 10'h009;
        mem[473] = 10'h27e;
        mem[474] = 10'h150;
        mem[475] = 10'h0b6;
        mem[476] = 10'h348;
        mem[477] = 10'h3f6;
        mem[478] = 10'h047;
        mem[479] = 10'h155;
        mem[480] = 10'h212;
        mem[481] = 10'h137;
        mem[482] = 10'h116;
        mem[483] = 10'h2fa;
        mem[484] = 10'h067;
        mem[485] = 10'h222;
        mem[486] = 10'h3c3;
        mem[487] = 10'h118;
        mem[488] = 10'h192;
        mem[489] = 10'h362;
        mem[490] = 10'h12d;
        mem[491] = 10'h361;
        mem[492] = 10'h3d0;
        mem[493] = 10'h2e7;
        mem[494] = 10'h338;
        mem[495] = 10'h285;
        mem[496] = 10'h0ce;
        mem[497] = 10'h27d;
        mem[498] = 10'h02a;
        mem[499] = 10'h122;
        mem[500] = 10'h2ea;
        mem[501] = 10'h316;
        mem[502] = 10'h16c;
        mem[503] = 10'h0ea;
        mem[504] = 10'h0dd;
        mem[505] = 10'h369;
        mem[506] = 10'h2d2;
        mem[507] = 10'h2c2;
        mem[508] = 10'h3da;
        mem[509] = 10'h295;
        mem[510] = 10'h180;
        mem[511] = 10'h21a;
        mem[512] = 10'h351;
        mem[513] = 10'h0be;
        mem[514] = 10'h041;
        mem[515] = 10'h3e5;
        mem[516] = 10'h13a;
        mem[517] = 10'h213;
        mem[518] = 10'h124;
        mem[519] = 10'h06a;
        mem[520] = 10'h278;
        mem[521] = 10'h04a;
        mem[522] = 10'h28b;
        mem[523] = 10'h117;
        mem[524] = 10'h319;
        mem[525] = 10'h023;
        mem[526] = 10'h162;
        mem[527] = 10'h3de;
        mem[528] = 10'h372;
        mem[529] = 10'h1da;
        mem[530] = 10'h120;
        mem[531] = 10'h0de;
        mem[532] = 10'h1bd;
        mem[533] = 10'h2f8;
        mem[534] = 10'h221;
        mem[535] = 10'h148;
        mem[536] = 10'h078;
        mem[537] = 10'h380;
        mem[538] = 10'h197;
        mem[539] = 10'h296;
        mem[540] = 10'h013;
        mem[541] = 10'h3ac;
        mem[542] = 10'h3f2;
        mem[543] = 10'h01d;
        mem[544] = 10'h22a;
        mem[545] = 10'h054;
        mem[546] = 10'h0f5;
        mem[547] = 10'h0bd;
        mem[548] = 10'h3e8;
        mem[549] = 10'h085;
        mem[550] = 10'h272;
        mem[551] = 10'h0e7;
        mem[552] = 10'h144;
        mem[553] = 10'h26f;
        mem[554] = 10'h391;
        mem[555] = 10'h113;
        mem[556] = 10'h3d5;
        mem[557] = 10'h1f3;
        mem[558] = 10'h3ee;
        mem[559] = 10'h38a;
        mem[560] = 10'h326;
        mem[561] = 10'h18e;
        mem[562] = 10'h0ca;
        mem[563] = 10'h226;
        mem[564] = 10'h236;
        mem[565] = 10'h1b0;
        mem[566] = 10'h119;
        mem[567] = 10'h2cf;
        mem[568] = 10'h19c;
        mem[569] = 10'h1dd;
        mem[570] = 10'h0d9;
        mem[571] = 10'h359;
        mem[572] = 10'h1cb;
        mem[573] = 10'h10d;
        mem[574] = 10'h16b;
        mem[575] = 10'h312;
        mem[576] = 10'h193;
        mem[577] = 10'h13e;
        mem[578] = 10'h11e;
        mem[579] = 10'h0ec;
        mem[580] = 10'h147;
        mem[581] = 10'h207;
        mem[582] = 10'h104;
        mem[583] = 10'h23a;
        mem[584] = 10'h166;
        mem[585] = 10'h289;
        mem[586] = 10'h07f;
        mem[587] = 10'h1e4;
        mem[588] = 10'h0b0;
        mem[589] = 10'h33e;
        mem[590] = 10'h175;
        mem[591] = 10'h10f;
        mem[592] = 10'h010;
        mem[593] = 10'h220;
        mem[594] = 10'h397;
        mem[595] = 10'h18c;
        mem[596] = 10'h294;
        mem[597] = 10'h145;
        mem[598] = 10'h014;
        mem[599] = 10'h2db;
        mem[600] = 10'h12a;
        mem[601] = 10'h099;
        mem[602] = 10'h129;
        mem[603] = 10'h389;
        mem[604] = 10'h282;
        mem[605] = 10'h195;
        mem[606] = 10'h1a3;
        mem[607] = 10'h268;
        mem[608] = 10'h320;
        mem[609] = 10'h0b4;
        mem[610] = 10'h3dd;
        mem[611] = 10'h1a9;
        mem[612] = 10'h005;
        mem[613] = 10'h339;
        mem[614] = 10'h241;
        mem[615] = 10'h1b6;
        mem[616] = 10'h2e9;
        mem[617] = 10'h363;
        mem[618] = 10'h21f;
        mem[619] = 10'h0c7;
        mem[620] = 10'h10a;
        mem[621] = 10'h250;
        mem[622] = 10'h1f1;
        mem[623] = 10'h073;
        mem[624] = 10'h28e;
        mem[625] = 10'h112;
        mem[626] = 10'h1cd;
        mem[627] = 10'h281;
        mem[628] = 10'h3d7;
        mem[629] = 10'h0eb;
        mem[630] = 10'h39a;
        mem[631] = 10'h108;
        mem[632] = 10'h09d;
        mem[633] = 10'h30f;
        mem[634] = 10'h105;
        mem[635] = 10'h2f4;
        mem[636] = 10'h1ad;
        mem[637] = 10'h17c;
        mem[638] = 10'h01a;
        mem[639] = 10'h0da;
        mem[640] = 10'h364;
        mem[641] = 10'h2a2;
        mem[642] = 10'h1dc;
        mem[643] = 10'h1b3;
        mem[644] = 10'h090;
        mem[645] = 10'h132;
        mem[646] = 10'h3e6;
        mem[647] = 10'h06c;
        mem[648] = 10'h1c4;
        mem[649] = 10'h15e;
        mem[650] = 10'h25d;
        mem[651] = 10'h0e9;
        mem[652] = 10'h0d5;
        mem[653] = 10'h0f1;
        mem[654] = 10'h043;
        mem[655] = 10'h083;
        mem[656] = 10'h21b;
        mem[657] = 10'h029;
        mem[658] = 10'h237;
        mem[659] = 10'h356;
        mem[660] = 10'h301;
        mem[661] = 10'h153;
        mem[662] = 10'h3fb;
        mem[663] = 10'h070;
        mem[664] = 10'h34f;
        mem[665] = 10'h23e;
        mem[666] = 10'h02f;
        mem[667] = 10'h32d;
        mem[668] = 10'h265;
        mem[669] = 10'h290;
        mem[670] = 10'h172;
        mem[671] = 10'h3e7;
        mem[672] = 10'h097;
        mem[673] = 10'h2d7;
        mem[674] = 10'h140;
        mem[675] = 10'h089;
        mem[676] = 10'h0fd;
        mem[677] = 10'h37e;
        mem[678] = 10'h3c5;
        mem[679] = 10'h2be;
        mem[680] = 10'h18f;
        mem[681] = 10'h1d8;
        mem[682] = 10'h164;
        mem[683] = 10'h038;
        mem[684] = 10'h20a;
        mem[685] = 10'h39b;
        mem[686] = 10'h22c;
        mem[687] = 10'h2c8;
        mem[688] = 10'h0fb;
        mem[689] = 10'h016;
        mem[690] = 10'h2fd;
        mem[691] = 10'h321;
        mem[692] = 10'h1d5;
        mem[693] = 10'h26c;
        mem[694] = 10'h218;
        mem[695] = 10'h292;
        mem[696] = 10'h354;
        mem[697] = 10'h29f;
        mem[698] = 10'h11a;
        mem[699] = 10'h0f2;
        mem[700] = 10'h26e;
        mem[701] = 10'h30a;
        mem[702] = 10'h2ce;
        mem[703] = 10'h185;
        mem[704] = 10'h165;
        mem[705] = 10'h2d1;
        mem[706] = 10'h08b;
        mem[707] = 10'h245;
        mem[708] = 10'h2ef;
        mem[709] = 10'h38b;
        mem[710] = 10'h28f;
        mem[711] = 10'h2d8;
        mem[712] = 10'h358;
        mem[713] = 10'h26b;
        mem[714] = 10'h3a7;
        mem[715] = 10'h0f3;
        mem[716] = 10'h3c8;
        mem[717] = 10'h086;
        mem[718] = 10'h1fc;
        mem[719] = 10'h224;
        mem[720] = 10'h1be;
        mem[721] = 10'h254;
        mem[722] = 10'h3c2;
        mem[723] = 10'h1bb;
        mem[724] = 10'h0bb;
        mem[725] = 10'h14e;
        mem[726] = 10'h398;
        mem[727] = 10'h06e;
        mem[728] = 10'h329;
        mem[729] = 10'h1de;
        mem[730] = 10'h1fd;
        mem[731] = 10'h19a;
        mem[732] = 10'h37b;
        mem[733] = 10'h229;
        mem[734] = 10'h058;
        mem[735] = 10'h399;
        mem[736] = 10'h303;
        mem[737] = 10'h123;
        mem[738] = 10'h03c;
        mem[739] = 10'h36c;
        mem[740] = 10'h201;
        mem[741] = 10'h395;
        mem[742] = 10'h0b7;
        mem[743] = 10'h028;
        mem[744] = 10'h05f;
        mem[745] = 10'h23c;
        mem[746] = 10'h0ef;
        mem[747] = 10'h0fa;
        mem[748] = 10'h3d4;
        mem[749] = 10'h3fc;
        mem[750] = 10'h05e;
        mem[751] = 10'h253;
        mem[752] = 10'h1d4;
        mem[753] = 10'h3a5;
        mem[754] = 10'h024;
        mem[755] = 10'h05a;
        mem[756] = 10'h127;
        mem[757] = 10'h161;
        mem[758] = 10'h1c5;
        mem[759] = 10'h035;
        mem[760] = 10'h27c;
        mem[761] = 10'h02b;
        mem[762] = 10'h1c6;
        mem[763] = 10'h152;
        mem[764] = 10'h018;
        mem[765] = 10'h3e9;
        mem[766] = 10'h146;
        mem[767] = 10'h2a7;
        mem[768] = 10'h048;
        mem[769] = 10'h219;
        mem[770] = 10'h37a;
        mem[771] = 10'h15d;
        mem[772] = 10'h388;
        mem[773] = 10'h293;
        mem[774] = 10'h0a8;
        mem[775] = 10'h333;
        mem[776] = 10'h3bf;
        mem[777] = 10'h020;
        mem[778] = 10'h199;
        mem[779] = 10'h12e;
        mem[780] = 10'h0d8;
        mem[781] = 10'h17e;
        mem[782] = 10'h3b2;
        mem[783] = 10'h2c4;
        mem[784] = 10'h196;
        mem[785] = 10'h366;
        mem[786] = 10'h3c1;
        mem[787] = 10'h05b;
        mem[788] = 10'h280;
        mem[789] = 10'h00b;
        mem[790] = 10'h02e;
        mem[791] = 10'h111;
        mem[792] = 10'h238;
        mem[793] = 10'h0a6;
        mem[794] = 10'h3bd;
        mem[795] = 10'h0a4;
        mem[796] = 10'h328;
        mem[797] = 10'h331;
        mem[798] = 10'h14d;
        mem[799] = 10'h15f;
        mem[800] = 10'h22d;
        mem[801] = 10'h2cc;
        mem[802] = 10'h353;
        mem[803] = 10'h2a1;
        mem[804] = 10'h1c8;
        mem[805] = 10'h286;
        mem[806] = 10'h313;
        mem[807] = 10'h08f;
        mem[808] = 10'h2f0;
        mem[809] = 10'h2a6;
        mem[810] = 10'h298;
        mem[811] = 10'h35e;
        mem[812] = 10'h271;
        mem[813] = 10'h381;
        mem[814] = 10'h171;
        mem[815] = 10'h2d0;
        mem[816] = 10'h3e1;
        mem[817] = 10'h0a9;
        mem[818] = 10'h38f;
        mem[819] = 10'h0d0;
        mem[820] = 10'h3ad;
        mem[821] = 10'h181;
        mem[822] = 10'h1df;
        mem[823] = 10'h346;
        mem[824] = 10'h098;
        mem[825] = 10'h1b5;
        mem[826] = 10'h374;
        mem[827] = 10'h30e;
        mem[828] = 10'h35c;
        mem[829] = 10'h13b;
        mem[830] = 10'h283;
        mem[831] = 10'h0d4;
        mem[832] = 10'h12c;
        mem[833] = 10'h1cc;
        mem[834] = 10'h2e6;
        mem[835] = 10'h0db;
        mem[836] = 10'h1ce;
        mem[837] = 10'h069;
        mem[838] = 10'h1ec;
        mem[839] = 10'h3b0;
        mem[840] = 10'h32b;
        mem[841] = 10'h34a;
        mem[842] = 10'h36d;
        mem[843] = 10'h05c;
        mem[844] = 10'h2da;
        mem[845] = 10'h183;
        mem[846] = 10'h230;
        mem[847] = 10'h3eb;
        mem[848] = 10'h121;
        mem[849] = 10'h15c;
        mem[850] = 10'h1d2;
        mem[851] = 10'h004;
        mem[852] = 10'h125;
        mem[853] = 10'h077;
        mem[854] = 10'h1b8;
        mem[855] = 10'h030;
        mem[856] = 10'h31c;
        mem[857] = 10'h2d5;
        mem[858] = 10'h1e6;
        mem[859] = 10'h39d;
        mem[860] = 10'h3d8;
        mem[861] = 10'h00a;
        mem[862] = 10'h142;
        mem[863] = 10'h209;
        mem[864] = 10'h09e;
        mem[865] = 10'h106;
        mem[866] = 10'h033;
        mem[867] = 10'h09b;
        mem[868] = 10'h1e9;
        mem[869] = 10'h215;
        mem[870] = 10'h1b9;
        mem[871] = 10'h367;
        mem[872] = 10'h159;
        mem[873] = 10'h32a;
        mem[874] = 10'h188;
        mem[875] = 10'h335;
        mem[876] = 10'h093;
        mem[877] = 10'h04b;
        mem[878] = 10'h3b5;
        mem[879] = 10'h2b1;
        mem[880] = 10'h35f;
        mem[881] = 10'h088;
        mem[882] = 10'h025;
        mem[883] = 10'h3b3;
        mem[884] = 10'h1fb;
        mem[885] = 10'h2cb;
        mem[886] = 10'h307;
        mem[887] = 10'h039;
        mem[888] = 10'h342;
        mem[889] = 10'h102;
        mem[890] = 10'h053;
        mem[891] = 10'h29a;
        mem[892] = 10'h276;
        mem[893] = 10'h3df;
        mem[894] = 10'h28a;
        mem[895] = 10'h288;
        mem[896] = 10'h341;
        mem[897] = 10'h042;
        mem[898] = 10'h360;
        mem[899] = 10'h1e8;
        mem[900] = 10'h071;
        mem[901] = 10'h3ff;
        mem[902] = 10'h01f;
        mem[903] = 10'h2f7;
        mem[904] = 10'h16d;
        mem[905] = 10'h00c;
        mem[906] = 10'h003;
        mem[907] = 10'h0c2;
        mem[908] = 10'h252;
        mem[909] = 10'h3f3;
        mem[910] = 10'h012;
        mem[911] = 10'h274;
        mem[912] = 10'h0ad;
        mem[913] = 10'h050;
        mem[914] = 10'h24d;
        mem[915] = 10'h1a1;
        mem[916] = 10'h141;
        mem[917] = 10'h154;
        mem[918] = 10'h344;
        mem[919] = 10'h2b7;
        mem[920] = 10'h136;
        mem[921] = 10'h27f;
        mem[922] = 10'h128;
        mem[923] = 10'h055;
        mem[924] = 10'h176;
        mem[925] = 10'h2b9;
        mem[926] = 10'h382;
        mem[927] = 10'h0e2;
        mem[928] = 10'h25b;
        mem[929] = 10'h25f;
        mem[930] = 10'h103;
        mem[931] = 10'h056;
        mem[932] = 10'h327;
        mem[933] = 10'h08a;
        mem[934] = 10'h1ea;
        mem[935] = 10'h310;
        mem[936] = 10'h081;
        mem[937] = 10'h0c1;
        mem[938] = 10'h244;
        mem[939] = 10'h2df;
        mem[940] = 10'h2d9;
        mem[941] = 10'h1f2;
        mem[942] = 10'h149;
        mem[943] = 10'h110;
        mem[944] = 10'h22e;
        mem[945] = 10'h034;
        mem[946] = 10'h080;
        mem[947] = 10'h0e3;
        mem[948] = 10'h18a;
        mem[949] = 10'h2ba;
        mem[950] = 10'h20b;
        mem[951] = 10'h357;
        mem[952] = 10'h2dc;
        mem[953] = 10'h28d;
        mem[954] = 10'h29d;
        mem[955] = 10'h16f;
        mem[956] = 10'h037;
        mem[957] = 10'h0a0;
        mem[958] = 10'h3f9;
        mem[959] = 10'h2e0;
        mem[960] = 10'h38e;
        mem[961] = 10'h091;
        mem[962] = 10'h13d;
        mem[963] = 10'h2f9;
        mem[964] = 10'h1a2;
        mem[965] = 10'h2c3;
        mem[966] = 10'h1a4;
        mem[967] = 10'h34e;
        mem[968] = 10'h002;
        mem[969] = 10'h0a5;
        mem[970] = 10'h163;
        mem[971] = 10'h062;
        mem[972] = 10'h1bf;
        mem[973] = 10'h14c;
        mem[974] = 10'h21c;
        mem[975] = 10'h0b9;
        mem[976] = 10'h107;
        mem[977] = 10'h06b;
        mem[978] = 10'h051;
        mem[979] = 10'h0c9;
        mem[980] = 10'h072;
        mem[981] = 10'h3f0;
        mem[982] = 10'h04c;
        mem[983] = 10'h3dc;
        mem[984] = 10'h065;
        mem[985] = 10'h2fc;
        mem[986] = 10'h3f8;
        mem[987] = 10'h14a;
        mem[988] = 10'h173;
        mem[989] = 10'h36b;
        mem[990] = 10'h31d;
        mem[991] = 10'h370;
        mem[992] = 10'h2f6;
        mem[993] = 10'h322;
        mem[994] = 10'h24b;
        mem[995] = 10'h206;
        mem[996] = 10'h0ff;
        mem[997] = 10'h157;
        mem[998] = 10'h170;
        mem[999] = 10'h373;
        mem[1000] = 10'h255;
        mem[1001] = 10'h115;
        mem[1002] = 10'h0e6;
        mem[1003] = 10'h32c;
        mem[1004] = 10'h1d7;
        mem[1005] = 10'h3b4;
        mem[1006] = 10'h0b2;
        mem[1007] = 10'h349;
        mem[1008] = 10'h3d3;
        mem[1009] = 10'h2ca;
        mem[1010] = 10'h34c;
        mem[1011] = 10'h2ed;
        mem[1012] = 10'h087;
        mem[1013] = 10'h304;
        mem[1014] = 10'h34b;
        mem[1015] = 10'h19e;
        mem[1016] = 10'h2b8;
        mem[1017] = 10'h0aa;
        mem[1018] = 10'h3a8;
        mem[1019] = 10'h03f;
        mem[1020] = 10'h291;
        mem[1021] = 10'h0d2;
        mem[1022] = 10'h036;
        mem[1023] = 10'h045;
    end
endmodule

module encrypt_4sbox_large6(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h105;
        mem[1] = 10'h2d5;
        mem[2] = 10'h3b8;
        mem[3] = 10'h383;
        mem[4] = 10'h27b;
        mem[5] = 10'h17f;
        mem[6] = 10'h0db;
        mem[7] = 10'h1ad;
        mem[8] = 10'h221;
        mem[9] = 10'h23f;
        mem[10] = 10'h042;
        mem[11] = 10'h089;
        mem[12] = 10'h1d5;
        mem[13] = 10'h0a3;
        mem[14] = 10'h3e5;
        mem[15] = 10'h14f;
        mem[16] = 10'h17d;
        mem[17] = 10'h125;
        mem[18] = 10'h1ba;
        mem[19] = 10'h040;
        mem[20] = 10'h33c;
        mem[21] = 10'h18b;
        mem[22] = 10'h3e9;
        mem[23] = 10'h118;
        mem[24] = 10'h011;
        mem[25] = 10'h21a;
        mem[26] = 10'h21f;
        mem[27] = 10'h29f;
        mem[28] = 10'h35e;
        mem[29] = 10'h3f6;
        mem[30] = 10'h063;
        mem[31] = 10'h0f2;
        mem[32] = 10'h30d;
        mem[33] = 10'h327;
        mem[34] = 10'h095;
        mem[35] = 10'h2bb;
        mem[36] = 10'h27d;
        mem[37] = 10'h020;
        mem[38] = 10'h052;
        mem[39] = 10'h22f;
        mem[40] = 10'h01b;
        mem[41] = 10'h0f0;
        mem[42] = 10'h2e0;
        mem[43] = 10'h312;
        mem[44] = 10'h250;
        mem[45] = 10'h2f0;
        mem[46] = 10'h171;
        mem[47] = 10'h3b5;
        mem[48] = 10'h05d;
        mem[49] = 10'h2d4;
        mem[50] = 10'h116;
        mem[51] = 10'h209;
        mem[52] = 10'h10a;
        mem[53] = 10'h235;
        mem[54] = 10'h2c8;
        mem[55] = 10'h1db;
        mem[56] = 10'h177;
        mem[57] = 10'h3fe;
        mem[58] = 10'h245;
        mem[59] = 10'h39f;
        mem[60] = 10'h02e;
        mem[61] = 10'h01a;
        mem[62] = 10'h2c7;
        mem[63] = 10'h01d;
        mem[64] = 10'h0eb;
        mem[65] = 10'h058;
        mem[66] = 10'h2a6;
        mem[67] = 10'h216;
        mem[68] = 10'h1b8;
        mem[69] = 10'h28e;
        mem[70] = 10'h121;
        mem[71] = 10'h28c;
        mem[72] = 10'h2db;
        mem[73] = 10'h1f9;
        mem[74] = 10'h2c2;
        mem[75] = 10'h38a;
        mem[76] = 10'h3d7;
        mem[77] = 10'h397;
        mem[78] = 10'h231;
        mem[79] = 10'h146;
        mem[80] = 10'h263;
        mem[81] = 10'h14a;
        mem[82] = 10'h199;
        mem[83] = 10'h251;
        mem[84] = 10'h0e1;
        mem[85] = 10'h1cf;
        mem[86] = 10'h24d;
        mem[87] = 10'h069;
        mem[88] = 10'h2cd;
        mem[89] = 10'h22e;
        mem[90] = 10'h1c4;
        mem[91] = 10'h2b8;
        mem[92] = 10'h19d;
        mem[93] = 10'h396;
        mem[94] = 10'h306;
        mem[95] = 10'h3c8;
        mem[96] = 10'h3c2;
        mem[97] = 10'h354;
        mem[98] = 10'h04d;
        mem[99] = 10'h1d4;
        mem[100] = 10'h28b;
        mem[101] = 10'h3ae;
        mem[102] = 10'h3c3;
        mem[103] = 10'h02f;
        mem[104] = 10'h1c3;
        mem[105] = 10'h359;
        mem[106] = 10'h2a7;
        mem[107] = 10'h060;
        mem[108] = 10'h094;
        mem[109] = 10'h127;
        mem[110] = 10'h154;
        mem[111] = 10'h176;
        mem[112] = 10'h281;
        mem[113] = 10'h02c;
        mem[114] = 10'h275;
        mem[115] = 10'h3c6;
        mem[116] = 10'h13c;
        mem[117] = 10'h376;
        mem[118] = 10'h0e7;
        mem[119] = 10'h344;
        mem[120] = 10'h025;
        mem[121] = 10'h0ce;
        mem[122] = 10'h11a;
        mem[123] = 10'h2e6;
        mem[124] = 10'h04c;
        mem[125] = 10'h336;
        mem[126] = 10'h096;
        mem[127] = 10'h236;
        mem[128] = 10'h38c;
        mem[129] = 10'h38e;
        mem[130] = 10'h07e;
        mem[131] = 10'h320;
        mem[132] = 10'h1e4;
        mem[133] = 10'h17b;
        mem[134] = 10'h375;
        mem[135] = 10'h11c;
        mem[136] = 10'h093;
        mem[137] = 10'h355;
        mem[138] = 10'h0e8;
        mem[139] = 10'h37d;
        mem[140] = 10'h2d2;
        mem[141] = 10'h13d;
        mem[142] = 10'h1c8;
        mem[143] = 10'h157;
        mem[144] = 10'h01c;
        mem[145] = 10'h009;
        mem[146] = 10'h341;
        mem[147] = 10'h3b4;
        mem[148] = 10'h1bc;
        mem[149] = 10'h29c;
        mem[150] = 10'h331;
        mem[151] = 10'h223;
        mem[152] = 10'h08c;
        mem[153] = 10'h3a9;
        mem[154] = 10'h212;
        mem[155] = 10'h192;
        mem[156] = 10'h126;
        mem[157] = 10'h039;
        mem[158] = 10'h1a3;
        mem[159] = 10'h180;
        mem[160] = 10'h34b;
        mem[161] = 10'h11e;
        mem[162] = 10'h1f1;
        mem[163] = 10'h2af;
        mem[164] = 10'h2be;
        mem[165] = 10'h1a5;
        mem[166] = 10'h178;
        mem[167] = 10'h003;
        mem[168] = 10'h3a4;
        mem[169] = 10'h30e;
        mem[170] = 10'h284;
        mem[171] = 10'h047;
        mem[172] = 10'h22a;
        mem[173] = 10'h3e6;
        mem[174] = 10'h357;
        mem[175] = 10'h0b3;
        mem[176] = 10'h2e2;
        mem[177] = 10'h218;
        mem[178] = 10'h1a2;
        mem[179] = 10'h2d9;
        mem[180] = 10'h198;
        mem[181] = 10'h117;
        mem[182] = 10'h3eb;
        mem[183] = 10'h252;
        mem[184] = 10'h377;
        mem[185] = 10'h1ae;
        mem[186] = 10'h22c;
        mem[187] = 10'h202;
        mem[188] = 10'h1f2;
        mem[189] = 10'h10e;
        mem[190] = 10'h005;
        mem[191] = 10'h1fb;
        mem[192] = 10'h267;
        mem[193] = 10'h1e5;
        mem[194] = 10'h0ed;
        mem[195] = 10'h33e;
        mem[196] = 10'h3da;
        mem[197] = 10'h0f6;
        mem[198] = 10'h072;
        mem[199] = 10'h352;
        mem[200] = 10'h124;
        mem[201] = 10'h2e9;
        mem[202] = 10'h32b;
        mem[203] = 10'h0ca;
        mem[204] = 10'h2bd;
        mem[205] = 10'h3a6;
        mem[206] = 10'h3af;
        mem[207] = 10'h06f;
        mem[208] = 10'h0b8;
        mem[209] = 10'h21c;
        mem[210] = 10'h150;
        mem[211] = 10'h3bd;
        mem[212] = 10'h0c5;
        mem[213] = 10'h391;
        mem[214] = 10'h140;
        mem[215] = 10'h373;
        mem[216] = 10'h3a3;
        mem[217] = 10'h269;
        mem[218] = 10'h2a8;
        mem[219] = 10'h16c;
        mem[220] = 10'h0a9;
        mem[221] = 10'h0a1;
        mem[222] = 10'h0bf;
        mem[223] = 10'h12a;
        mem[224] = 10'h385;
        mem[225] = 10'h1f7;
        mem[226] = 10'h1c0;
        mem[227] = 10'h276;
        mem[228] = 10'h2ee;
        mem[229] = 10'h0b7;
        mem[230] = 10'h298;
        mem[231] = 10'h0ef;
        mem[232] = 10'h274;
        mem[233] = 10'h064;
        mem[234] = 10'h0dc;
        mem[235] = 10'h00d;
        mem[236] = 10'h128;
        mem[237] = 10'h381;
        mem[238] = 10'h3db;
        mem[239] = 10'h25a;
        mem[240] = 10'h2a4;
        mem[241] = 10'h12c;
        mem[242] = 10'h074;
        mem[243] = 10'h3ec;
        mem[244] = 10'h101;
        mem[245] = 10'h3fd;
        mem[246] = 10'h23c;
        mem[247] = 10'h195;
        mem[248] = 10'h0ac;
        mem[249] = 10'h3c1;
        mem[250] = 10'h17e;
        mem[251] = 10'h00e;
        mem[252] = 10'h271;
        mem[253] = 10'h1d6;
        mem[254] = 10'h05e;
        mem[255] = 10'h270;
        mem[256] = 10'h01f;
        mem[257] = 10'h0d5;
        mem[258] = 10'h0ff;
        mem[259] = 10'h043;
        mem[260] = 10'h048;
        mem[261] = 10'h120;
        mem[262] = 10'h09b;
        mem[263] = 10'h16e;
        mem[264] = 10'h211;
        mem[265] = 10'h3d8;
        mem[266] = 10'h254;
        mem[267] = 10'h238;
        mem[268] = 10'h141;
        mem[269] = 10'h332;
        mem[270] = 10'h384;
        mem[271] = 10'h08e;
        mem[272] = 10'h335;
        mem[273] = 10'h315;
        mem[274] = 10'h3d5;
        mem[275] = 10'h1c5;
        mem[276] = 10'h1c7;
        mem[277] = 10'h0cd;
        mem[278] = 10'h309;
        mem[279] = 10'h36f;
        mem[280] = 10'h3ac;
        mem[281] = 10'h00f;
        mem[282] = 10'h1aa;
        mem[283] = 10'h350;
        mem[284] = 10'h25e;
        mem[285] = 10'h2d7;
        mem[286] = 10'h110;
        mem[287] = 10'h188;
        mem[288] = 10'h260;
        mem[289] = 10'h019;
        mem[290] = 10'h104;
        mem[291] = 10'h3ef;
        mem[292] = 10'h2e8;
        mem[293] = 10'h079;
        mem[294] = 10'h34d;
        mem[295] = 10'h225;
        mem[296] = 10'h081;
        mem[297] = 10'h2ae;
        mem[298] = 10'h03f;
        mem[299] = 10'h380;
        mem[300] = 10'h1c9;
        mem[301] = 10'h000;
        mem[302] = 10'h1eb;
        mem[303] = 10'h001;
        mem[304] = 10'h015;
        mem[305] = 10'h307;
        mem[306] = 10'h389;
        mem[307] = 10'h3f7;
        mem[308] = 10'h076;
        mem[309] = 10'h205;
        mem[310] = 10'h37c;
        mem[311] = 10'h246;
        mem[312] = 10'h02b;
        mem[313] = 10'h394;
        mem[314] = 10'h179;
        mem[315] = 10'h186;
        mem[316] = 10'h129;
        mem[317] = 10'h2b0;
        mem[318] = 10'h3ba;
        mem[319] = 10'h2cc;
        mem[320] = 10'h155;
        mem[321] = 10'h09c;
        mem[322] = 10'h322;
        mem[323] = 10'h214;
        mem[324] = 10'h3a1;
        mem[325] = 10'h39d;
        mem[326] = 10'h2d0;
        mem[327] = 10'h1ec;
        mem[328] = 10'h0f7;
        mem[329] = 10'h030;
        mem[330] = 10'h1a9;
        mem[331] = 10'h2aa;
        mem[332] = 10'h25b;
        mem[333] = 10'h061;
        mem[334] = 10'h326;
        mem[335] = 10'h1f5;
        mem[336] = 10'h36e;
        mem[337] = 10'h356;
        mem[338] = 10'h256;
        mem[339] = 10'h207;
        mem[340] = 10'h3a7;
        mem[341] = 10'h220;
        mem[342] = 10'h3cd;
        mem[343] = 10'h091;
        mem[344] = 10'h1f0;
        mem[345] = 10'h143;
        mem[346] = 10'h172;
        mem[347] = 10'h32a;
        mem[348] = 10'h185;
        mem[349] = 10'h1d3;
        mem[350] = 10'h15f;
        mem[351] = 10'h1bd;
        mem[352] = 10'h1cc;
        mem[353] = 10'h277;
        mem[354] = 10'h0a4;
        mem[355] = 10'h227;
        mem[356] = 10'h37f;
        mem[357] = 10'h2b3;
        mem[358] = 10'h398;
        mem[359] = 10'h3d3;
        mem[360] = 10'h0e9;
        mem[361] = 10'h0c9;
        mem[362] = 10'h145;
        mem[363] = 10'h20b;
        mem[364] = 10'h343;
        mem[365] = 10'h149;
        mem[366] = 10'h1fa;
        mem[367] = 10'h1d1;
        mem[368] = 10'h3c7;
        mem[369] = 10'h06d;
        mem[370] = 10'h25f;
        mem[371] = 10'h229;
        mem[372] = 10'h0c1;
        mem[373] = 10'h258;
        mem[374] = 10'h365;
        mem[375] = 10'h0b6;
        mem[376] = 10'h2ec;
        mem[377] = 10'h15e;
        mem[378] = 10'h282;
        mem[379] = 10'h337;
        mem[380] = 10'h0aa;
        mem[381] = 10'h388;
        mem[382] = 10'h29e;
        mem[383] = 10'h20f;
        mem[384] = 10'h2b4;
        mem[385] = 10'h2f2;
        mem[386] = 10'h1cd;
        mem[387] = 10'h12b;
        mem[388] = 10'h2ba;
        mem[389] = 10'h296;
        mem[390] = 10'h374;
        mem[391] = 10'h390;
        mem[392] = 10'h173;
        mem[393] = 10'h2e3;
        mem[394] = 10'h106;
        mem[395] = 10'h316;
        mem[396] = 10'h334;
        mem[397] = 10'h3cb;
        mem[398] = 10'h1d0;
        mem[399] = 10'h0d0;
        mem[400] = 10'h082;
        mem[401] = 10'h2b2;
        mem[402] = 10'h0de;
        mem[403] = 10'h1a0;
        mem[404] = 10'h289;
        mem[405] = 10'h05b;
        mem[406] = 10'h1b5;
        mem[407] = 10'h392;
        mem[408] = 10'h10c;
        mem[409] = 10'h23d;
        mem[410] = 10'h090;
        mem[411] = 10'h35f;
        mem[412] = 10'h13a;
        mem[413] = 10'h305;
        mem[414] = 10'h0c7;
        mem[415] = 10'h136;
        mem[416] = 10'h39c;
        mem[417] = 10'h370;
        mem[418] = 10'h1d8;
        mem[419] = 10'h1a1;
        mem[420] = 10'h097;
        mem[421] = 10'h313;
        mem[422] = 10'h166;
        mem[423] = 10'h314;
        mem[424] = 10'h273;
        mem[425] = 10'h3fa;
        mem[426] = 10'h24e;
        mem[427] = 10'h18f;
        mem[428] = 10'h2fb;
        mem[429] = 10'h2f6;
        mem[430] = 10'h3d2;
        mem[431] = 10'h193;
        mem[432] = 10'h2eb;
        mem[433] = 10'h33f;
        mem[434] = 10'h0be;
        mem[435] = 10'h31b;
        mem[436] = 10'h26e;
        mem[437] = 10'h37e;
        mem[438] = 10'h18d;
        mem[439] = 10'h19b;
        mem[440] = 10'h36c;
        mem[441] = 10'h20e;
        mem[442] = 10'h295;
        mem[443] = 10'h02a;
        mem[444] = 10'h280;
        mem[445] = 10'h0f1;
        mem[446] = 10'h2a5;
        mem[447] = 10'h0c3;
        mem[448] = 10'h36b;
        mem[449] = 10'h3e4;
        mem[450] = 10'h37b;
        mem[451] = 10'h018;
        mem[452] = 10'h15c;
        mem[453] = 10'h2c5;
        mem[454] = 10'h299;
        mem[455] = 10'h272;
        mem[456] = 10'h0d6;
        mem[457] = 10'h0e2;
        mem[458] = 10'h16d;
        mem[459] = 10'h22d;
        mem[460] = 10'h028;
        mem[461] = 10'h09a;
        mem[462] = 10'h107;
        mem[463] = 10'h0c2;
        mem[464] = 10'h302;
        mem[465] = 10'h0b1;
        mem[466] = 10'h168;
        mem[467] = 10'h0ae;
        mem[468] = 10'h04a;
        mem[469] = 10'h2f4;
        mem[470] = 10'h163;
        mem[471] = 10'h0c8;
        mem[472] = 10'h31d;
        mem[473] = 10'h1c1;
        mem[474] = 10'h2d6;
        mem[475] = 10'h059;
        mem[476] = 10'h15b;
        mem[477] = 10'h0c6;
        mem[478] = 10'h2b6;
        mem[479] = 10'h197;
        mem[480] = 10'h03c;
        mem[481] = 10'h07c;
        mem[482] = 10'h240;
        mem[483] = 10'h26b;
        mem[484] = 10'h1ca;
        mem[485] = 10'h24c;
        mem[486] = 10'h054;
        mem[487] = 10'h1d2;
        mem[488] = 10'h098;
        mem[489] = 10'h213;
        mem[490] = 10'h08f;
        mem[491] = 10'h1e1;
        mem[492] = 10'h14c;
        mem[493] = 10'h215;
        mem[494] = 10'h30a;
        mem[495] = 10'h0b5;
        mem[496] = 10'h2d1;
        mem[497] = 10'h055;
        mem[498] = 10'h2f5;
        mem[499] = 10'h0c4;
        mem[500] = 10'h290;
        mem[501] = 10'h3c9;
        mem[502] = 10'h050;
        mem[503] = 10'h0e6;
        mem[504] = 10'h1fe;
        mem[505] = 10'h234;
        mem[506] = 10'h2bc;
        mem[507] = 10'h0d7;
        mem[508] = 10'h3ea;
        mem[509] = 10'h1bb;
        mem[510] = 10'h1e3;
        mem[511] = 10'h21b;
        mem[512] = 10'h008;
        mem[513] = 10'h137;
        mem[514] = 10'h17c;
        mem[515] = 10'h349;
        mem[516] = 10'h1b0;
        mem[517] = 10'h0bd;
        mem[518] = 10'h05a;
        mem[519] = 10'h0e0;
        mem[520] = 10'h037;
        mem[521] = 10'h0ec;
        mem[522] = 10'h3ab;
        mem[523] = 10'h1b9;
        mem[524] = 10'h28a;
        mem[525] = 10'h333;
        mem[526] = 10'h18e;
        mem[527] = 10'h268;
        mem[528] = 10'h024;
        mem[529] = 10'h387;
        mem[530] = 10'h078;
        mem[531] = 10'h0f8;
        mem[532] = 10'h294;
        mem[533] = 10'h23a;
        mem[534] = 10'h0ab;
        mem[535] = 10'h2b9;
        mem[536] = 10'h1e7;
        mem[537] = 10'h2ed;
        mem[538] = 10'h0f3;
        mem[539] = 10'h367;
        mem[540] = 10'h3dd;
        mem[541] = 10'h06b;
        mem[542] = 10'h2e7;
        mem[543] = 10'h080;
        mem[544] = 10'h2c6;
        mem[545] = 10'h051;
        mem[546] = 10'h070;
        mem[547] = 10'h113;
        mem[548] = 10'h03e;
        mem[549] = 10'h288;
        mem[550] = 10'h2fd;
        mem[551] = 10'h39a;
        mem[552] = 10'h099;
        mem[553] = 10'h181;
        mem[554] = 10'h162;
        mem[555] = 10'h0fa;
        mem[556] = 10'h23b;
        mem[557] = 10'h0ee;
        mem[558] = 10'h36a;
        mem[559] = 10'h368;
        mem[560] = 10'h2a0;
        mem[561] = 10'h190;
        mem[562] = 10'h0d8;
        mem[563] = 10'h07d;
        mem[564] = 10'h0fd;
        mem[565] = 10'h395;
        mem[566] = 10'h14d;
        mem[567] = 10'h28d;
        mem[568] = 10'h0a7;
        mem[569] = 10'h1ef;
        mem[570] = 10'h3d4;
        mem[571] = 10'h175;
        mem[572] = 10'h264;
        mem[573] = 10'h27c;
        mem[574] = 10'h3ad;
        mem[575] = 10'h293;
        mem[576] = 10'h353;
        mem[577] = 10'h39b;
        mem[578] = 10'h297;
        mem[579] = 10'h364;
        mem[580] = 10'h347;
        mem[581] = 10'h3bb;
        mem[582] = 10'h33a;
        mem[583] = 10'h13e;
        mem[584] = 10'h26d;
        mem[585] = 10'h217;
        mem[586] = 10'h1f4;
        mem[587] = 10'h0b0;
        mem[588] = 10'h3e0;
        mem[589] = 10'h012;
        mem[590] = 10'h2de;
        mem[591] = 10'h24f;
        mem[592] = 10'h369;
        mem[593] = 10'h386;
        mem[594] = 10'h1a8;
        mem[595] = 10'h242;
        mem[596] = 10'h1a6;
        mem[597] = 10'h2d8;
        mem[598] = 10'h100;
        mem[599] = 10'h0e3;
        mem[600] = 10'h0dd;
        mem[601] = 10'h362;
        mem[602] = 10'h31f;
        mem[603] = 10'h021;
        mem[604] = 10'h0d4;
        mem[605] = 10'h036;
        mem[606] = 10'h378;
        mem[607] = 10'h3f2;
        mem[608] = 10'h38d;
        mem[609] = 10'h261;
        mem[610] = 10'h027;
        mem[611] = 10'h21d;
        mem[612] = 10'h1d7;
        mem[613] = 10'h133;
        mem[614] = 10'h0fc;
        mem[615] = 10'h3f4;
        mem[616] = 10'h138;
        mem[617] = 10'h3a0;
        mem[618] = 10'h148;
        mem[619] = 10'h32e;
        mem[620] = 10'h346;
        mem[621] = 10'h2ab;
        mem[622] = 10'h3b2;
        mem[623] = 10'h3b7;
        mem[624] = 10'h329;
        mem[625] = 10'h3f0;
        mem[626] = 10'h1b4;
        mem[627] = 10'h085;
        mem[628] = 10'h2f7;
        mem[629] = 10'h19f;
        mem[630] = 10'h3b6;
        mem[631] = 10'h0f5;
        mem[632] = 10'h3e1;
        mem[633] = 10'h187;
        mem[634] = 10'h04e;
        mem[635] = 10'h210;
        mem[636] = 10'h067;
        mem[637] = 10'h366;
        mem[638] = 10'h3e8;
        mem[639] = 10'h170;
        mem[640] = 10'h318;
        mem[641] = 10'h10f;
        mem[642] = 10'h2c0;
        mem[643] = 10'h0f9;
        mem[644] = 10'h35d;
        mem[645] = 10'h27a;
        mem[646] = 10'h371;
        mem[647] = 10'h244;
        mem[648] = 10'h1b3;
        mem[649] = 10'h248;
        mem[650] = 10'h3cf;
        mem[651] = 10'h07f;
        mem[652] = 10'h132;
        mem[653] = 10'h233;
        mem[654] = 10'h071;
        mem[655] = 10'h32f;
        mem[656] = 10'h123;
        mem[657] = 10'h158;
        mem[658] = 10'h03a;
        mem[659] = 10'h372;
        mem[660] = 10'h32d;
        mem[661] = 10'h08a;
        mem[662] = 10'h30c;
        mem[663] = 10'h249;
        mem[664] = 10'h1ff;
        mem[665] = 10'h1cb;
        mem[666] = 10'h0ea;
        mem[667] = 10'h108;
        mem[668] = 10'h2e4;
        mem[669] = 10'h2c9;
        mem[670] = 10'h34e;
        mem[671] = 10'h3ff;
        mem[672] = 10'h0fb;
        mem[673] = 10'h27f;
        mem[674] = 10'h339;
        mem[675] = 10'h382;
        mem[676] = 10'h12e;
        mem[677] = 10'h262;
        mem[678] = 10'h363;
        mem[679] = 10'h11b;
        mem[680] = 10'h144;
        mem[681] = 10'h35b;
        mem[682] = 10'h2dc;
        mem[683] = 10'h09d;
        mem[684] = 10'h301;
        mem[685] = 10'h303;
        mem[686] = 10'h2cb;
        mem[687] = 10'h230;
        mem[688] = 10'h075;
        mem[689] = 10'h109;
        mem[690] = 10'h33d;
        mem[691] = 10'h08b;
        mem[692] = 10'h183;
        mem[693] = 10'h204;
        mem[694] = 10'h134;
        mem[695] = 10'h0bb;
        mem[696] = 10'h399;
        mem[697] = 10'h0b9;
        mem[698] = 10'h19e;
        mem[699] = 10'h1e9;
        mem[700] = 10'h09f;
        mem[701] = 10'h3e3;
        mem[702] = 10'h04b;
        mem[703] = 10'h345;
        mem[704] = 10'h3c4;
        mem[705] = 10'h35a;
        mem[706] = 10'h1de;
        mem[707] = 10'h013;
        mem[708] = 10'h2f3;
        mem[709] = 10'h1da;
        mem[710] = 10'h21e;
        mem[711] = 10'h029;
        mem[712] = 10'h3fb;
        mem[713] = 10'h0a6;
        mem[714] = 10'h3f5;
        mem[715] = 10'h286;
        mem[716] = 10'h3c0;
        mem[717] = 10'h2f9;
        mem[718] = 10'h304;
        mem[719] = 10'h1b6;
        mem[720] = 10'h135;
        mem[721] = 10'h19c;
        mem[722] = 10'h161;
        mem[723] = 10'h1c6;
        mem[724] = 10'h330;
        mem[725] = 10'h39e;
        mem[726] = 10'h285;
        mem[727] = 10'h0a5;
        mem[728] = 10'h08d;
        mem[729] = 10'h26f;
        mem[730] = 10'h310;
        mem[731] = 10'h2bf;
        mem[732] = 10'h073;
        mem[733] = 10'h004;
        mem[734] = 10'h0cf;
        mem[735] = 10'h1b2;
        mem[736] = 10'h3dc;
        mem[737] = 10'h328;
        mem[738] = 10'h31c;
        mem[739] = 10'h253;
        mem[740] = 10'h0f4;
        mem[741] = 10'h278;
        mem[742] = 10'h3bc;
        mem[743] = 10'h26c;
        mem[744] = 10'h0d1;
        mem[745] = 10'h142;
        mem[746] = 10'h088;
        mem[747] = 10'h07b;
        mem[748] = 10'h0c0;
        mem[749] = 10'h0a2;
        mem[750] = 10'h07a;
        mem[751] = 10'h182;
        mem[752] = 10'h15a;
        mem[753] = 10'h010;
        mem[754] = 10'h3b1;
        mem[755] = 10'h29a;
        mem[756] = 10'h1dc;
        mem[757] = 10'h152;
        mem[758] = 10'h10d;
        mem[759] = 10'h2a9;
        mem[760] = 10'h26a;
        mem[761] = 10'h2d3;
        mem[762] = 10'h10b;
        mem[763] = 10'h131;
        mem[764] = 10'h00c;
        mem[765] = 10'h02d;
        mem[766] = 10'h0a8;
        mem[767] = 10'h3b9;
        mem[768] = 10'h3f9;
        mem[769] = 10'h114;
        mem[770] = 10'h1fc;
        mem[771] = 10'h38f;
        mem[772] = 10'h20d;
        mem[773] = 10'h393;
        mem[774] = 10'h044;
        mem[775] = 10'h1e0;
        mem[776] = 10'h1af;
        mem[777] = 10'h122;
        mem[778] = 10'h1e6;
        mem[779] = 10'h15d;
        mem[780] = 10'h1f6;
        mem[781] = 10'h006;
        mem[782] = 10'h3cc;
        mem[783] = 10'h196;
        mem[784] = 10'h053;
        mem[785] = 10'h30f;
        mem[786] = 10'h045;
        mem[787] = 10'h2ce;
        mem[788] = 10'h16b;
        mem[789] = 10'h2dd;
        mem[790] = 10'h1ee;
        mem[791] = 10'h228;
        mem[792] = 10'h1ac;
        mem[793] = 10'h28f;
        mem[794] = 10'h201;
        mem[795] = 10'h3ee;
        mem[796] = 10'h017;
        mem[797] = 10'h17a;
        mem[798] = 10'h007;
        mem[799] = 10'h33b;
        mem[800] = 10'h086;
        mem[801] = 10'h1f8;
        mem[802] = 10'h16a;
        mem[803] = 10'h29b;
        mem[804] = 10'h0af;
        mem[805] = 10'h062;
        mem[806] = 10'h27e;
        mem[807] = 10'h3bf;
        mem[808] = 10'h292;
        mem[809] = 10'h184;
        mem[810] = 10'h169;
        mem[811] = 10'h014;
        mem[812] = 10'h1b7;
        mem[813] = 10'h200;
        mem[814] = 10'h3aa;
        mem[815] = 10'h283;
        mem[816] = 10'h1ed;
        mem[817] = 10'h156;
        mem[818] = 10'h0cc;
        mem[819] = 10'h226;
        mem[820] = 10'h041;
        mem[821] = 10'h119;
        mem[822] = 10'h2fa;
        mem[823] = 10'h3f3;
        mem[824] = 10'h317;
        mem[825] = 10'h1dd;
        mem[826] = 10'h3d1;
        mem[827] = 10'h379;
        mem[828] = 10'h083;
        mem[829] = 10'h3d6;
        mem[830] = 10'h241;
        mem[831] = 10'h3a5;
        mem[832] = 10'h13b;
        mem[833] = 10'h324;
        mem[834] = 10'h01e;
        mem[835] = 10'h189;
        mem[836] = 10'h2da;
        mem[837] = 10'h342;
        mem[838] = 10'h102;
        mem[839] = 10'h20a;
        mem[840] = 10'h11d;
        mem[841] = 10'h300;
        mem[842] = 10'h3ca;
        mem[843] = 10'h2a1;
        mem[844] = 10'h167;
        mem[845] = 10'h3be;
        mem[846] = 10'h321;
        mem[847] = 10'h159;
        mem[848] = 10'h29d;
        mem[849] = 10'h3ce;
        mem[850] = 10'h077;
        mem[851] = 10'h092;
        mem[852] = 10'h255;
        mem[853] = 10'h139;
        mem[854] = 10'h348;
        mem[855] = 10'h084;
        mem[856] = 10'h115;
        mem[857] = 10'h11f;
        mem[858] = 10'h2c1;
        mem[859] = 10'h2ac;
        mem[860] = 10'h2b7;
        mem[861] = 10'h066;
        mem[862] = 10'h338;
        mem[863] = 10'h3a2;
        mem[864] = 10'h023;
        mem[865] = 10'h243;
        mem[866] = 10'h0e5;
        mem[867] = 10'h32c;
        mem[868] = 10'h37a;
        mem[869] = 10'h0a0;
        mem[870] = 10'h291;
        mem[871] = 10'h206;
        mem[872] = 10'h3e2;
        mem[873] = 10'h3f8;
        mem[874] = 10'h03b;
        mem[875] = 10'h1a7;
        mem[876] = 10'h239;
        mem[877] = 10'h2e1;
        mem[878] = 10'h34a;
        mem[879] = 10'h032;
        mem[880] = 10'h1bf;
        mem[881] = 10'h2a3;
        mem[882] = 10'h1d9;
        mem[883] = 10'h237;
        mem[884] = 10'h03d;
        mem[885] = 10'h3e7;
        mem[886] = 10'h00a;
        mem[887] = 10'h0ba;
        mem[888] = 10'h1b1;
        mem[889] = 10'h0cb;
        mem[890] = 10'h265;
        mem[891] = 10'h1be;
        mem[892] = 10'h034;
        mem[893] = 10'h20c;
        mem[894] = 10'h1e2;
        mem[895] = 10'h222;
        mem[896] = 10'h153;
        mem[897] = 10'h038;
        mem[898] = 10'h002;
        mem[899] = 10'h112;
        mem[900] = 10'h3c5;
        mem[901] = 10'h30b;
        mem[902] = 10'h164;
        mem[903] = 10'h0e4;
        mem[904] = 10'h319;
        mem[905] = 10'h0ad;
        mem[906] = 10'h2a2;
        mem[907] = 10'h34c;
        mem[908] = 10'h24b;
        mem[909] = 10'h1ab;
        mem[910] = 10'h1ea;
        mem[911] = 10'h016;
        mem[912] = 10'h360;
        mem[913] = 10'h087;
        mem[914] = 10'h358;
        mem[915] = 10'h25c;
        mem[916] = 10'h0d2;
        mem[917] = 10'h3d0;
        mem[918] = 10'h0b2;
        mem[919] = 10'h1ce;
        mem[920] = 10'h022;
        mem[921] = 10'h2e5;
        mem[922] = 10'h18c;
        mem[923] = 10'h031;
        mem[924] = 10'h1fd;
        mem[925] = 10'h0d9;
        mem[926] = 10'h06c;
        mem[927] = 10'h130;
        mem[928] = 10'h068;
        mem[929] = 10'h09e;
        mem[930] = 10'h3a8;
        mem[931] = 10'h0b4;
        mem[932] = 10'h2f1;
        mem[933] = 10'h194;
        mem[934] = 10'h340;
        mem[935] = 10'h2c3;
        mem[936] = 10'h36d;
        mem[937] = 10'h035;
        mem[938] = 10'h247;
        mem[939] = 10'h34f;
        mem[940] = 10'h311;
        mem[941] = 10'h23e;
        mem[942] = 10'h06e;
        mem[943] = 10'h219;
        mem[944] = 10'h3fc;
        mem[945] = 10'h208;
        mem[946] = 10'h05c;
        mem[947] = 10'h2b1;
        mem[948] = 10'h325;
        mem[949] = 10'h103;
        mem[950] = 10'h165;
        mem[951] = 10'h259;
        mem[952] = 10'h13f;
        mem[953] = 10'h224;
        mem[954] = 10'h31a;
        mem[955] = 10'h06a;
        mem[956] = 10'h0fe;
        mem[957] = 10'h12d;
        mem[958] = 10'h308;
        mem[959] = 10'h12f;
        mem[960] = 10'h25d;
        mem[961] = 10'h3b3;
        mem[962] = 10'h232;
        mem[963] = 10'h2cf;
        mem[964] = 10'h323;
        mem[965] = 10'h3d9;
        mem[966] = 10'h2c4;
        mem[967] = 10'h361;
        mem[968] = 10'h065;
        mem[969] = 10'h0bc;
        mem[970] = 10'h1a4;
        mem[971] = 10'h3ed;
        mem[972] = 10'h3f1;
        mem[973] = 10'h266;
        mem[974] = 10'h026;
        mem[975] = 10'h3df;
        mem[976] = 10'h057;
        mem[977] = 10'h1e8;
        mem[978] = 10'h18a;
        mem[979] = 10'h2ca;
        mem[980] = 10'h174;
        mem[981] = 10'h160;
        mem[982] = 10'h22b;
        mem[983] = 10'h191;
        mem[984] = 10'h2b5;
        mem[985] = 10'h351;
        mem[986] = 10'h31e;
        mem[987] = 10'h35c;
        mem[988] = 10'h033;
        mem[989] = 10'h00b;
        mem[990] = 10'h3b0;
        mem[991] = 10'h046;
        mem[992] = 10'h3de;
        mem[993] = 10'h056;
        mem[994] = 10'h111;
        mem[995] = 10'h05f;
        mem[996] = 10'h2fc;
        mem[997] = 10'h2ff;
        mem[998] = 10'h2f8;
        mem[999] = 10'h0df;
        mem[1000] = 10'h1df;
        mem[1001] = 10'h14e;
        mem[1002] = 10'h279;
        mem[1003] = 10'h151;
        mem[1004] = 10'h2ad;
        mem[1005] = 10'h2df;
        mem[1006] = 10'h04f;
        mem[1007] = 10'h2fe;
        mem[1008] = 10'h147;
        mem[1009] = 10'h287;
        mem[1010] = 10'h257;
        mem[1011] = 10'h14b;
        mem[1012] = 10'h38b;
        mem[1013] = 10'h1c2;
        mem[1014] = 10'h16f;
        mem[1015] = 10'h2ea;
        mem[1016] = 10'h203;
        mem[1017] = 10'h1f3;
        mem[1018] = 10'h2ef;
        mem[1019] = 10'h0d3;
        mem[1020] = 10'h0da;
        mem[1021] = 10'h049;
        mem[1022] = 10'h19a;
        mem[1023] = 10'h24a;
    end
endmodule

module encrypt_4sbox_large7(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h17d;
        mem[1] = 10'h0d0;
        mem[2] = 10'h1cc;
        mem[3] = 10'h1fd;
        mem[4] = 10'h0a0;
        mem[5] = 10'h28f;
        mem[6] = 10'h32d;
        mem[7] = 10'h3fe;
        mem[8] = 10'h0f2;
        mem[9] = 10'h142;
        mem[10] = 10'h3d8;
        mem[11] = 10'h2ea;
        mem[12] = 10'h141;
        mem[13] = 10'h27b;
        mem[14] = 10'h0c0;
        mem[15] = 10'h2df;
        mem[16] = 10'h13c;
        mem[17] = 10'h393;
        mem[18] = 10'h08e;
        mem[19] = 10'h024;
        mem[20] = 10'h24c;
        mem[21] = 10'h272;
        mem[22] = 10'h1d1;
        mem[23] = 10'h39f;
        mem[24] = 10'h2ab;
        mem[25] = 10'h339;
        mem[26] = 10'h175;
        mem[27] = 10'h081;
        mem[28] = 10'h3d5;
        mem[29] = 10'h157;
        mem[30] = 10'h086;
        mem[31] = 10'h28a;
        mem[32] = 10'h3d2;
        mem[33] = 10'h255;
        mem[34] = 10'h1b4;
        mem[35] = 10'h2d2;
        mem[36] = 10'h034;
        mem[37] = 10'h256;
        mem[38] = 10'h317;
        mem[39] = 10'h3ab;
        mem[40] = 10'h1d3;
        mem[41] = 10'h163;
        mem[42] = 10'h0d5;
        mem[43] = 10'h16e;
        mem[44] = 10'h05e;
        mem[45] = 10'h18a;
        mem[46] = 10'h3f9;
        mem[47] = 10'h209;
        mem[48] = 10'h2b2;
        mem[49] = 10'h080;
        mem[50] = 10'h051;
        mem[51] = 10'h3dc;
        mem[52] = 10'h287;
        mem[53] = 10'h130;
        mem[54] = 10'h00c;
        mem[55] = 10'h20c;
        mem[56] = 10'h3ba;
        mem[57] = 10'h3fc;
        mem[58] = 10'h1a0;
        mem[59] = 10'h05c;
        mem[60] = 10'h19b;
        mem[61] = 10'h25d;
        mem[62] = 10'h09c;
        mem[63] = 10'h0c1;
        mem[64] = 10'h12f;
        mem[65] = 10'h220;
        mem[66] = 10'h34e;
        mem[67] = 10'h216;
        mem[68] = 10'h1d8;
        mem[69] = 10'h0d9;
        mem[70] = 10'h3e6;
        mem[71] = 10'h36e;
        mem[72] = 10'h02a;
        mem[73] = 10'h003;
        mem[74] = 10'h109;
        mem[75] = 10'h22b;
        mem[76] = 10'h311;
        mem[77] = 10'h2f6;
        mem[78] = 10'h366;
        mem[79] = 10'h016;
        mem[80] = 10'h143;
        mem[81] = 10'h3fd;
        mem[82] = 10'h026;
        mem[83] = 10'h0f3;
        mem[84] = 10'h065;
        mem[85] = 10'h07f;
        mem[86] = 10'h147;
        mem[87] = 10'h1e1;
        mem[88] = 10'h100;
        mem[89] = 10'h171;
        mem[90] = 10'h35b;
        mem[91] = 10'h083;
        mem[92] = 10'h16c;
        mem[93] = 10'h07c;
        mem[94] = 10'h0a3;
        mem[95] = 10'h32e;
        mem[96] = 10'h3ca;
        mem[97] = 10'h0f1;
        mem[98] = 10'h164;
        mem[99] = 10'h129;
        mem[100] = 10'h225;
        mem[101] = 10'h153;
        mem[102] = 10'h36d;
        mem[103] = 10'h0e1;
        mem[104] = 10'h041;
        mem[105] = 10'h0c4;
        mem[106] = 10'h12b;
        mem[107] = 10'h18f;
        mem[108] = 10'h038;
        mem[109] = 10'h073;
        mem[110] = 10'h087;
        mem[111] = 10'h0af;
        mem[112] = 10'h2bc;
        mem[113] = 10'h07b;
        mem[114] = 10'h2aa;
        mem[115] = 10'h2ba;
        mem[116] = 10'h0df;
        mem[117] = 10'h296;
        mem[118] = 10'h24e;
        mem[119] = 10'h0ed;
        mem[120] = 10'h181;
        mem[121] = 10'h31a;
        mem[122] = 10'h33a;
        mem[123] = 10'h358;
        mem[124] = 10'h154;
        mem[125] = 10'h2ee;
        mem[126] = 10'h302;
        mem[127] = 10'h2e3;
        mem[128] = 10'h168;
        mem[129] = 10'h38d;
        mem[130] = 10'h1ad;
        mem[131] = 10'h1d5;
        mem[132] = 10'h152;
        mem[133] = 10'h11d;
        mem[134] = 10'h01f;
        mem[135] = 10'h353;
        mem[136] = 10'h1a1;
        mem[137] = 10'h11f;
        mem[138] = 10'h2a3;
        mem[139] = 10'h230;
        mem[140] = 10'h39b;
        mem[141] = 10'h0de;
        mem[142] = 10'h218;
        mem[143] = 10'h2b1;
        mem[144] = 10'h24b;
        mem[145] = 10'h0bf;
        mem[146] = 10'h294;
        mem[147] = 10'h3e2;
        mem[148] = 10'h099;
        mem[149] = 10'h115;
        mem[150] = 10'h30a;
        mem[151] = 10'h08d;
        mem[152] = 10'h261;
        mem[153] = 10'h3a8;
        mem[154] = 10'h0e4;
        mem[155] = 10'h2da;
        mem[156] = 10'h37e;
        mem[157] = 10'h2f1;
        mem[158] = 10'h258;
        mem[159] = 10'h3d1;
        mem[160] = 10'h1ba;
        mem[161] = 10'h1b0;
        mem[162] = 10'h1a9;
        mem[163] = 10'h161;
        mem[164] = 10'h1cb;
        mem[165] = 10'h1ff;
        mem[166] = 10'h31d;
        mem[167] = 10'h3fa;
        mem[168] = 10'h193;
        mem[169] = 10'h155;
        mem[170] = 10'h336;
        mem[171] = 10'h203;
        mem[172] = 10'h08c;
        mem[173] = 10'h098;
        mem[174] = 10'h177;
        mem[175] = 10'h34d;
        mem[176] = 10'h208;
        mem[177] = 10'h05b;
        mem[178] = 10'h330;
        mem[179] = 10'h3ac;
        mem[180] = 10'h02c;
        mem[181] = 10'h382;
        mem[182] = 10'h1cf;
        mem[183] = 10'h09b;
        mem[184] = 10'h013;
        mem[185] = 10'h328;
        mem[186] = 10'h361;
        mem[187] = 10'h38a;
        mem[188] = 10'h1c3;
        mem[189] = 10'h31c;
        mem[190] = 10'h29c;
        mem[191] = 10'h039;
        mem[192] = 10'h032;
        mem[193] = 10'h273;
        mem[194] = 10'h079;
        mem[195] = 10'h368;
        mem[196] = 10'h0f9;
        mem[197] = 10'h0e3;
        mem[198] = 10'h375;
        mem[199] = 10'h160;
        mem[200] = 10'h2cb;
        mem[201] = 10'h332;
        mem[202] = 10'h117;
        mem[203] = 10'h2dc;
        mem[204] = 10'h289;
        mem[205] = 10'h396;
        mem[206] = 10'h151;
        mem[207] = 10'h2d8;
        mem[208] = 10'h14b;
        mem[209] = 10'h30c;
        mem[210] = 10'h3f6;
        mem[211] = 10'h14f;
        mem[212] = 10'h06d;
        mem[213] = 10'h1ab;
        mem[214] = 10'h126;
        mem[215] = 10'h352;
        mem[216] = 10'h2f5;
        mem[217] = 10'h18b;
        mem[218] = 10'h1f8;
        mem[219] = 10'h190;
        mem[220] = 10'h1a5;
        mem[221] = 10'h07d;
        mem[222] = 10'h3df;
        mem[223] = 10'h0d3;
        mem[224] = 10'h263;
        mem[225] = 10'h3ce;
        mem[226] = 10'h377;
        mem[227] = 10'h124;
        mem[228] = 10'h245;
        mem[229] = 10'h194;
        mem[230] = 10'h315;
        mem[231] = 10'h1e3;
        mem[232] = 10'h223;
        mem[233] = 10'h379;
        mem[234] = 10'h188;
        mem[235] = 10'h1c0;
        mem[236] = 10'h1ed;
        mem[237] = 10'h0d8;
        mem[238] = 10'h351;
        mem[239] = 10'h2c4;
        mem[240] = 10'h090;
        mem[241] = 10'h0ba;
        mem[242] = 10'h3cc;
        mem[243] = 10'h269;
        mem[244] = 10'h105;
        mem[245] = 10'h3a1;
        mem[246] = 10'h133;
        mem[247] = 10'h1c6;
        mem[248] = 10'h13b;
        mem[249] = 10'h2f0;
        mem[250] = 10'h15a;
        mem[251] = 10'h023;
        mem[252] = 10'h36f;
        mem[253] = 10'h191;
        mem[254] = 10'h347;
        mem[255] = 10'h1ac;
        mem[256] = 10'h2ff;
        mem[257] = 10'h21c;
        mem[258] = 10'h227;
        mem[259] = 10'h01b;
        mem[260] = 10'h32b;
        mem[261] = 10'h2be;
        mem[262] = 10'h185;
        mem[263] = 10'h242;
        mem[264] = 10'h2ef;
        mem[265] = 10'h217;
        mem[266] = 10'h2b7;
        mem[267] = 10'h094;
        mem[268] = 10'h342;
        mem[269] = 10'h002;
        mem[270] = 10'h0a5;
        mem[271] = 10'h380;
        mem[272] = 10'h20e;
        mem[273] = 10'h2c9;
        mem[274] = 10'h3ad;
        mem[275] = 10'h0ee;
        mem[276] = 10'h2de;
        mem[277] = 10'h101;
        mem[278] = 10'h3a0;
        mem[279] = 10'h28c;
        mem[280] = 10'h096;
        mem[281] = 10'h0c7;
        mem[282] = 10'h048;
        mem[283] = 10'h06c;
        mem[284] = 10'h32f;
        mem[285] = 10'h355;
        mem[286] = 10'h314;
        mem[287] = 10'h310;
        mem[288] = 10'h265;
        mem[289] = 10'h20f;
        mem[290] = 10'h39c;
        mem[291] = 10'h20d;
        mem[292] = 10'h308;
        mem[293] = 10'h350;
        mem[294] = 10'h14c;
        mem[295] = 10'h0b5;
        mem[296] = 10'h1f3;
        mem[297] = 10'h089;
        mem[298] = 10'h0f0;
        mem[299] = 10'h138;
        mem[300] = 10'h3db;
        mem[301] = 10'h057;
        mem[302] = 10'h224;
        mem[303] = 10'h291;
        mem[304] = 10'h307;
        mem[305] = 10'h316;
        mem[306] = 10'h23f;
        mem[307] = 10'h3c8;
        mem[308] = 10'h39e;
        mem[309] = 10'h33d;
        mem[310] = 10'h3e5;
        mem[311] = 10'h159;
        mem[312] = 10'h0da;
        mem[313] = 10'h2ce;
        mem[314] = 10'h030;
        mem[315] = 10'h0a9;
        mem[316] = 10'h367;
        mem[317] = 10'h3cf;
        mem[318] = 10'h03a;
        mem[319] = 10'h278;
        mem[320] = 10'h006;
        mem[321] = 10'h06a;
        mem[322] = 10'h2fe;
        mem[323] = 10'h318;
        mem[324] = 10'h01c;
        mem[325] = 10'h025;
        mem[326] = 10'h3b9;
        mem[327] = 10'h288;
        mem[328] = 10'h0f4;
        mem[329] = 10'h2f4;
        mem[330] = 10'h00b;
        mem[331] = 10'h3da;
        mem[332] = 10'h3e4;
        mem[333] = 10'h3ff;
        mem[334] = 10'h166;
        mem[335] = 10'h12c;
        mem[336] = 10'h16d;
        mem[337] = 10'h173;
        mem[338] = 10'h1a3;
        mem[339] = 10'h30b;
        mem[340] = 10'h11c;
        mem[341] = 10'h240;
        mem[342] = 10'h01a;
        mem[343] = 10'h2b4;
        mem[344] = 10'h3a4;
        mem[345] = 10'h390;
        mem[346] = 10'h3c5;
        mem[347] = 10'h35e;
        mem[348] = 10'h077;
        mem[349] = 10'h2f7;
        mem[350] = 10'h274;
        mem[351] = 10'h211;
        mem[352] = 10'h1ee;
        mem[353] = 10'h144;
        mem[354] = 10'h2f3;
        mem[355] = 10'h0b9;
        mem[356] = 10'h276;
        mem[357] = 10'h386;
        mem[358] = 10'h07a;
        mem[359] = 10'h0cd;
        mem[360] = 10'h1f2;
        mem[361] = 10'h36c;
        mem[362] = 10'h2a8;
        mem[363] = 10'h1ec;
        mem[364] = 10'h058;
        mem[365] = 10'h3aa;
        mem[366] = 10'h075;
        mem[367] = 10'h200;
        mem[368] = 10'h248;
        mem[369] = 10'h0a8;
        mem[370] = 10'h365;
        mem[371] = 10'h1c2;
        mem[372] = 10'h114;
        mem[373] = 10'h162;
        mem[374] = 10'h1a4;
        mem[375] = 10'h2e9;
        mem[376] = 10'h1af;
        mem[377] = 10'h167;
        mem[378] = 10'h32a;
        mem[379] = 10'h035;
        mem[380] = 10'h2e5;
        mem[381] = 10'h3a9;
        mem[382] = 10'h3b7;
        mem[383] = 10'h1d2;
        mem[384] = 10'h360;
        mem[385] = 10'h2e0;
        mem[386] = 10'h183;
        mem[387] = 10'h088;
        mem[388] = 10'h14e;
        mem[389] = 10'h2a1;
        mem[390] = 10'h213;
        mem[391] = 10'h1aa;
        mem[392] = 10'h0ea;
        mem[393] = 10'h2fb;
        mem[394] = 10'h222;
        mem[395] = 10'h299;
        mem[396] = 10'h3b5;
        mem[397] = 10'h3a7;
        mem[398] = 10'h17b;
        mem[399] = 10'h1b1;
        mem[400] = 10'h362;
        mem[401] = 10'h37a;
        mem[402] = 10'h150;
        mem[403] = 10'h2fa;
        mem[404] = 10'h345;
        mem[405] = 10'h093;
        mem[406] = 10'h069;
        mem[407] = 10'h00a;
        mem[408] = 10'h322;
        mem[409] = 10'h313;
        mem[410] = 10'h04b;
        mem[411] = 10'h2dd;
        mem[412] = 10'h17a;
        mem[413] = 10'h0fe;
        mem[414] = 10'h33b;
        mem[415] = 10'h321;
        mem[416] = 10'h34c;
        mem[417] = 10'h2fd;
        mem[418] = 10'h028;
        mem[419] = 10'h16b;
        mem[420] = 10'h3b1;
        mem[421] = 10'h3b0;
        mem[422] = 10'h281;
        mem[423] = 10'h082;
        mem[424] = 10'h27f;
        mem[425] = 10'h2a2;
        mem[426] = 10'h37c;
        mem[427] = 10'h14d;
        mem[428] = 10'h195;
        mem[429] = 10'h264;
        mem[430] = 10'h054;
        mem[431] = 10'h26b;
        mem[432] = 10'h09f;
        mem[433] = 10'h19a;
        mem[434] = 10'h3bd;
        mem[435] = 10'h0e8;
        mem[436] = 10'h1f7;
        mem[437] = 10'h3c2;
        mem[438] = 10'h15d;
        mem[439] = 10'h019;
        mem[440] = 10'h2a4;
        mem[441] = 10'h2e2;
        mem[442] = 10'h04e;
        mem[443] = 10'h2ad;
        mem[444] = 10'h0a4;
        mem[445] = 10'h0db;
        mem[446] = 10'h325;
        mem[447] = 10'h135;
        mem[448] = 10'h27a;
        mem[449] = 10'h00d;
        mem[450] = 10'h306;
        mem[451] = 10'h285;
        mem[452] = 10'h13e;
        mem[453] = 10'h303;
        mem[454] = 10'h0cf;
        mem[455] = 10'h1f5;
        mem[456] = 10'h28b;
        mem[457] = 10'h280;
        mem[458] = 10'h1e0;
        mem[459] = 10'h03c;
        mem[460] = 10'h3f7;
        mem[461] = 10'h388;
        mem[462] = 10'h3c4;
        mem[463] = 10'h21a;
        mem[464] = 10'h1f1;
        mem[465] = 10'h049;
        mem[466] = 10'h29a;
        mem[467] = 10'h116;
        mem[468] = 10'h04c;
        mem[469] = 10'h06b;
        mem[470] = 10'h3b2;
        mem[471] = 10'h1b6;
        mem[472] = 10'h018;
        mem[473] = 10'h1da;
        mem[474] = 10'h28d;
        mem[475] = 10'h2c3;
        mem[476] = 10'h2e7;
        mem[477] = 10'h1a6;
        mem[478] = 10'h35d;
        mem[479] = 10'h38f;
        mem[480] = 10'h020;
        mem[481] = 10'h2cd;
        mem[482] = 10'h01d;
        mem[483] = 10'h15c;
        mem[484] = 10'h33f;
        mem[485] = 10'h25b;
        mem[486] = 10'h112;
        mem[487] = 10'h1e8;
        mem[488] = 10'h25a;
        mem[489] = 10'h2a6;
        mem[490] = 10'h1b8;
        mem[491] = 10'h34b;
        mem[492] = 10'h20a;
        mem[493] = 10'h1a7;
        mem[494] = 10'h22f;
        mem[495] = 10'h277;
        mem[496] = 10'h1ae;
        mem[497] = 10'h2d0;
        mem[498] = 10'h2c7;
        mem[499] = 10'h127;
        mem[500] = 10'h042;
        mem[501] = 10'h06e;
        mem[502] = 10'h128;
        mem[503] = 10'h2d5;
        mem[504] = 10'h12e;
        mem[505] = 10'h26e;
        mem[506] = 10'h13a;
        mem[507] = 10'h2e1;
        mem[508] = 10'h2d7;
        mem[509] = 10'h3f2;
        mem[510] = 10'h3ef;
        mem[511] = 10'h14a;
        mem[512] = 10'h0a2;
        mem[513] = 10'h0a1;
        mem[514] = 10'h305;
        mem[515] = 10'h0b8;
        mem[516] = 10'h0b7;
        mem[517] = 10'h219;
        mem[518] = 10'h2b5;
        mem[519] = 10'h338;
        mem[520] = 10'h346;
        mem[521] = 10'h1d9;
        mem[522] = 10'h2c2;
        mem[523] = 10'h0d2;
        mem[524] = 10'h23c;
        mem[525] = 10'h34f;
        mem[526] = 10'h207;
        mem[527] = 10'h085;
        mem[528] = 10'h0b4;
        mem[529] = 10'h0ca;
        mem[530] = 10'h071;
        mem[531] = 10'h010;
        mem[532] = 10'h097;
        mem[533] = 10'h229;
        mem[534] = 10'h3be;
        mem[535] = 10'h320;
        mem[536] = 10'h369;
        mem[537] = 10'h2bd;
        mem[538] = 10'h2a5;
        mem[539] = 10'h30d;
        mem[540] = 10'h10f;
        mem[541] = 10'h1ef;
        mem[542] = 10'h09d;
        mem[543] = 10'h247;
        mem[544] = 10'h275;
        mem[545] = 10'h045;
        mem[546] = 10'h012;
        mem[547] = 10'h148;
        mem[548] = 10'h20b;
        mem[549] = 10'h25f;
        mem[550] = 10'h16a;
        mem[551] = 10'h293;
        mem[552] = 10'h076;
        mem[553] = 10'h363;
        mem[554] = 10'h0eb;
        mem[555] = 10'h250;
        mem[556] = 10'h10e;
        mem[557] = 10'h033;
        mem[558] = 10'h3de;
        mem[559] = 10'h072;
        mem[560] = 10'h383;
        mem[561] = 10'h38b;
        mem[562] = 10'h2db;
        mem[563] = 10'h38e;
        mem[564] = 10'h02e;
        mem[565] = 10'h2a9;
        mem[566] = 10'h3e8;
        mem[567] = 10'h2ec;
        mem[568] = 10'h0fb;
        mem[569] = 10'h1e4;
        mem[570] = 10'h270;
        mem[571] = 10'h11a;
        mem[572] = 10'h23e;
        mem[573] = 10'h266;
        mem[574] = 10'h037;
        mem[575] = 10'h1c9;
        mem[576] = 10'h385;
        mem[577] = 10'h0e0;
        mem[578] = 10'h23d;
        mem[579] = 10'h286;
        mem[580] = 10'h074;
        mem[581] = 10'h119;
        mem[582] = 10'h2cc;
        mem[583] = 10'h1df;
        mem[584] = 10'h146;
        mem[585] = 10'h2d4;
        mem[586] = 10'h356;
        mem[587] = 10'h22c;
        mem[588] = 10'h047;
        mem[589] = 10'h331;
        mem[590] = 10'h254;
        mem[591] = 10'h1de;
        mem[592] = 10'h2d9;
        mem[593] = 10'h39d;
        mem[594] = 10'h2fc;
        mem[595] = 10'h18c;
        mem[596] = 10'h1b7;
        mem[597] = 10'h078;
        mem[598] = 10'h3cd;
        mem[599] = 10'h2b8;
        mem[600] = 10'h2f9;
        mem[601] = 10'h262;
        mem[602] = 10'h30f;
        mem[603] = 10'h1c5;
        mem[604] = 10'h205;
        mem[605] = 10'h1f9;
        mem[606] = 10'h1b5;
        mem[607] = 10'h1d6;
        mem[608] = 10'h060;
        mem[609] = 10'h21e;
        mem[610] = 10'h2b9;
        mem[611] = 10'h15b;
        mem[612] = 10'h27d;
        mem[613] = 10'h108;
        mem[614] = 10'h16f;
        mem[615] = 10'h050;
        mem[616] = 10'h0c8;
        mem[617] = 10'h169;
        mem[618] = 10'h397;
        mem[619] = 10'h297;
        mem[620] = 10'h004;
        mem[621] = 10'h0b1;
        mem[622] = 10'h206;
        mem[623] = 10'h0c6;
        mem[624] = 10'h13f;
        mem[625] = 10'h202;
        mem[626] = 10'h0f6;
        mem[627] = 10'h02f;
        mem[628] = 10'h0b2;
        mem[629] = 10'h3bf;
        mem[630] = 10'h235;
        mem[631] = 10'h267;
        mem[632] = 10'h172;
        mem[633] = 10'h29b;
        mem[634] = 10'h37f;
        mem[635] = 10'h131;
        mem[636] = 10'h246;
        mem[637] = 10'h1c8;
        mem[638] = 10'h10d;
        mem[639] = 10'h061;
        mem[640] = 10'h334;
        mem[641] = 10'h120;
        mem[642] = 10'h376;
        mem[643] = 10'h036;
        mem[644] = 10'h118;
        mem[645] = 10'h3ea;
        mem[646] = 10'h0b0;
        mem[647] = 10'h040;
        mem[648] = 10'h052;
        mem[649] = 10'h238;
        mem[650] = 10'h3f8;
        mem[651] = 10'h2af;
        mem[652] = 10'h139;
        mem[653] = 10'h29e;
        mem[654] = 10'h022;
        mem[655] = 10'h26a;
        mem[656] = 10'h0c2;
        mem[657] = 10'h03f;
        mem[658] = 10'h027;
        mem[659] = 10'h300;
        mem[660] = 10'h239;
        mem[661] = 10'h3c6;
        mem[662] = 10'h11e;
        mem[663] = 10'h24d;
        mem[664] = 10'h283;
        mem[665] = 10'h234;
        mem[666] = 10'h053;
        mem[667] = 10'h05d;
        mem[668] = 10'h22e;
        mem[669] = 10'h1e7;
        mem[670] = 10'h38c;
        mem[671] = 10'h1dc;
        mem[672] = 10'h237;
        mem[673] = 10'h0ec;
        mem[674] = 10'h08f;
        mem[675] = 10'h36b;
        mem[676] = 10'h106;
        mem[677] = 10'h103;
        mem[678] = 10'h387;
        mem[679] = 10'h309;
        mem[680] = 10'h2bb;
        mem[681] = 10'h0d7;
        mem[682] = 10'h295;
        mem[683] = 10'h189;
        mem[684] = 10'h19e;
        mem[685] = 10'h1f6;
        mem[686] = 10'h3c1;
        mem[687] = 10'h122;
        mem[688] = 10'h15e;
        mem[689] = 10'h3e0;
        mem[690] = 10'h3e1;
        mem[691] = 10'h1bc;
        mem[692] = 10'h1bb;
        mem[693] = 10'h3e3;
        mem[694] = 10'h3b8;
        mem[695] = 10'h0a6;
        mem[696] = 10'h374;
        mem[697] = 10'h02d;
        mem[698] = 10'h3af;
        mem[699] = 10'h125;
        mem[700] = 10'h066;
        mem[701] = 10'h29d;
        mem[702] = 10'h21d;
        mem[703] = 10'h12a;
        mem[704] = 10'h2f2;
        mem[705] = 10'h11b;
        mem[706] = 10'h3c7;
        mem[707] = 10'h31f;
        mem[708] = 10'h092;
        mem[709] = 10'h2ed;
        mem[710] = 10'h2ca;
        mem[711] = 10'h371;
        mem[712] = 10'h298;
        mem[713] = 10'h0e5;
        mem[714] = 10'h1a8;
        mem[715] = 10'h2c5;
        mem[716] = 10'h170;
        mem[717] = 10'h1d7;
        mem[718] = 10'h22d;
        mem[719] = 10'h1fe;
        mem[720] = 10'h0c3;
        mem[721] = 10'h1e5;
        mem[722] = 10'h3c3;
        mem[723] = 10'h134;
        mem[724] = 10'h2eb;
        mem[725] = 10'h381;
        mem[726] = 10'h21f;
        mem[727] = 10'h059;
        mem[728] = 10'h18d;
        mem[729] = 10'h043;
        mem[730] = 10'h228;
        mem[731] = 10'h1e9;
        mem[732] = 10'h0f5;
        mem[733] = 10'h2d1;
        mem[734] = 10'h35a;
        mem[735] = 10'h292;
        mem[736] = 10'h35f;
        mem[737] = 10'h0fc;
        mem[738] = 10'h327;
        mem[739] = 10'h26d;
        mem[740] = 10'h395;
        mem[741] = 10'h1d0;
        mem[742] = 10'h179;
        mem[743] = 10'h1bf;
        mem[744] = 10'h279;
        mem[745] = 10'h37d;
        mem[746] = 10'h132;
        mem[747] = 10'h1db;
        mem[748] = 10'h226;
        mem[749] = 10'h3e9;
        mem[750] = 10'h0d6;
        mem[751] = 10'h10a;
        mem[752] = 10'h09a;
        mem[753] = 10'h36a;
        mem[754] = 10'h319;
        mem[755] = 10'h28e;
        mem[756] = 10'h32c;
        mem[757] = 10'h337;
        mem[758] = 10'h3a6;
        mem[759] = 10'h196;
        mem[760] = 10'h199;
        mem[761] = 10'h354;
        mem[762] = 10'h31b;
        mem[763] = 10'h1dd;
        mem[764] = 10'h214;
        mem[765] = 10'h1e2;
        mem[766] = 10'h27c;
        mem[767] = 10'h136;
        mem[768] = 10'h22a;
        mem[769] = 10'h145;
        mem[770] = 10'h001;
        mem[771] = 10'h1be;
        mem[772] = 10'h2b0;
        mem[773] = 10'h243;
        mem[774] = 10'h253;
        mem[775] = 10'h1c4;
        mem[776] = 10'h23a;
        mem[777] = 10'h3c9;
        mem[778] = 10'h0dc;
        mem[779] = 10'h3a2;
        mem[780] = 10'h0dd;
        mem[781] = 10'h1ce;
        mem[782] = 10'h0ac;
        mem[783] = 10'h2c6;
        mem[784] = 10'h1b3;
        mem[785] = 10'h378;
        mem[786] = 10'h341;
        mem[787] = 10'h392;
        mem[788] = 10'h370;
        mem[789] = 10'h290;
        mem[790] = 10'h0fa;
        mem[791] = 10'h33e;
        mem[792] = 10'h0bd;
        mem[793] = 10'h156;
        mem[794] = 10'h2a7;
        mem[795] = 10'h27e;
        mem[796] = 10'h384;
        mem[797] = 10'h091;
        mem[798] = 10'h201;
        mem[799] = 10'h2f8;
        mem[800] = 10'h3bb;
        mem[801] = 10'h1fb;
        mem[802] = 10'h233;
        mem[803] = 10'h3d4;
        mem[804] = 10'h12d;
        mem[805] = 10'h21b;
        mem[806] = 10'h359;
        mem[807] = 10'h3f0;
        mem[808] = 10'h326;
        mem[809] = 10'h260;
        mem[810] = 10'h029;
        mem[811] = 10'h110;
        mem[812] = 10'h137;
        mem[813] = 10'h3ae;
        mem[814] = 10'h34a;
        mem[815] = 10'h187;
        mem[816] = 10'h05f;
        mem[817] = 10'h1f4;
        mem[818] = 10'h064;
        mem[819] = 10'h257;
        mem[820] = 10'h340;
        mem[821] = 10'h24a;
        mem[822] = 10'h249;
        mem[823] = 10'h212;
        mem[824] = 10'h215;
        mem[825] = 10'h3d9;
        mem[826] = 10'h17e;
        mem[827] = 10'h271;
        mem[828] = 10'h241;
        mem[829] = 10'h084;
        mem[830] = 10'h00e;
        mem[831] = 10'h07e;
        mem[832] = 10'h1bd;
        mem[833] = 10'h3d0;
        mem[834] = 10'h3f1;
        mem[835] = 10'h1a2;
        mem[836] = 10'h357;
        mem[837] = 10'h3dd;
        mem[838] = 10'h3ed;
        mem[839] = 10'h25c;
        mem[840] = 10'h04a;
        mem[841] = 10'h349;
        mem[842] = 10'h0fd;
        mem[843] = 10'h111;
        mem[844] = 10'h2e4;
        mem[845] = 10'h0e6;
        mem[846] = 10'h391;
        mem[847] = 10'h24f;
        mem[848] = 10'h0c5;
        mem[849] = 10'h2c0;
        mem[850] = 10'h008;
        mem[851] = 10'h372;
        mem[852] = 10'h1ca;
        mem[853] = 10'h3a5;
        mem[854] = 10'h1ea;
        mem[855] = 10'h0e7;
        mem[856] = 10'h0e9;
        mem[857] = 10'h09e;
        mem[858] = 10'h1b9;
        mem[859] = 10'h123;
        mem[860] = 10'h2ae;
        mem[861] = 10'h282;
        mem[862] = 10'h389;
        mem[863] = 10'h0cb;
        mem[864] = 10'h3eb;
        mem[865] = 10'h343;
        mem[866] = 10'h29f;
        mem[867] = 10'h121;
        mem[868] = 10'h165;
        mem[869] = 10'h0d4;
        mem[870] = 10'h015;
        mem[871] = 10'h0bc;
        mem[872] = 10'h18e;
        mem[873] = 10'h2b6;
        mem[874] = 10'h33c;
        mem[875] = 10'h04d;
        mem[876] = 10'h3ec;
        mem[877] = 10'h13d;
        mem[878] = 10'h301;
        mem[879] = 10'h03b;
        mem[880] = 10'h2ac;
        mem[881] = 10'h0f7;
        mem[882] = 10'h197;
        mem[883] = 10'h005;
        mem[884] = 10'h014;
        mem[885] = 10'h0f8;
        mem[886] = 10'h335;
        mem[887] = 10'h23b;
        mem[888] = 10'h232;
        mem[889] = 10'h15f;
        mem[890] = 10'h324;
        mem[891] = 10'h3b3;
        mem[892] = 10'h364;
        mem[893] = 10'h244;
        mem[894] = 10'h186;
        mem[895] = 10'h0ff;
        mem[896] = 10'h329;
        mem[897] = 10'h070;
        mem[898] = 10'h10c;
        mem[899] = 10'h398;
        mem[900] = 10'h210;
        mem[901] = 10'h176;
        mem[902] = 10'h021;
        mem[903] = 10'h158;
        mem[904] = 10'h2e6;
        mem[905] = 10'h174;
        mem[906] = 10'h26c;
        mem[907] = 10'h02b;
        mem[908] = 10'h05a;
        mem[909] = 10'h1cd;
        mem[910] = 10'h35c;
        mem[911] = 10'h3e7;
        mem[912] = 10'h0a7;
        mem[913] = 10'h19d;
        mem[914] = 10'h3cb;
        mem[915] = 10'h031;
        mem[916] = 10'h2d3;
        mem[917] = 10'h3f4;
        mem[918] = 10'h104;
        mem[919] = 10'h252;
        mem[920] = 10'h3c0;
        mem[921] = 10'h062;
        mem[922] = 10'h178;
        mem[923] = 10'h30e;
        mem[924] = 10'h0ae;
        mem[925] = 10'h1fa;
        mem[926] = 10'h3d7;
        mem[927] = 10'h17c;
        mem[928] = 10'h0ce;
        mem[929] = 10'h1c1;
        mem[930] = 10'h102;
        mem[931] = 10'h2c1;
        mem[932] = 10'h1b2;
        mem[933] = 10'h31e;
        mem[934] = 10'h0cc;
        mem[935] = 10'h068;
        mem[936] = 10'h1c7;
        mem[937] = 10'h0b6;
        mem[938] = 10'h046;
        mem[939] = 10'h007;
        mem[940] = 10'h348;
        mem[941] = 10'h2cf;
        mem[942] = 10'h182;
        mem[943] = 10'h3d6;
        mem[944] = 10'h236;
        mem[945] = 10'h067;
        mem[946] = 10'h198;
        mem[947] = 10'h056;
        mem[948] = 10'h0b3;
        mem[949] = 10'h1f0;
        mem[950] = 10'h3bc;
        mem[951] = 10'h2a0;
        mem[952] = 10'h0bb;
        mem[953] = 10'h3f5;
        mem[954] = 10'h0e2;
        mem[955] = 10'h0ad;
        mem[956] = 10'h25e;
        mem[957] = 10'h3f3;
        mem[958] = 10'h231;
        mem[959] = 10'h0ef;
        mem[960] = 10'h08a;
        mem[961] = 10'h044;
        mem[962] = 10'h140;
        mem[963] = 10'h19c;
        mem[964] = 10'h3b6;
        mem[965] = 10'h333;
        mem[966] = 10'h26f;
        mem[967] = 10'h2c8;
        mem[968] = 10'h0be;
        mem[969] = 10'h009;
        mem[970] = 10'h107;
        mem[971] = 10'h17f;
        mem[972] = 10'h01e;
        mem[973] = 10'h2e8;
        mem[974] = 10'h3fb;
        mem[975] = 10'h394;
        mem[976] = 10'h3ee;
        mem[977] = 10'h0d1;
        mem[978] = 10'h284;
        mem[979] = 10'h259;
        mem[980] = 10'h2bf;
        mem[981] = 10'h06f;
        mem[982] = 10'h323;
        mem[983] = 10'h19f;
        mem[984] = 10'h04f;
        mem[985] = 10'h063;
        mem[986] = 10'h0c9;
        mem[987] = 10'h149;
        mem[988] = 10'h0aa;
        mem[989] = 10'h10b;
        mem[990] = 10'h268;
        mem[991] = 10'h095;
        mem[992] = 10'h344;
        mem[993] = 10'h1e6;
        mem[994] = 10'h184;
        mem[995] = 10'h2b3;
        mem[996] = 10'h251;
        mem[997] = 10'h3b4;
        mem[998] = 10'h1fc;
        mem[999] = 10'h192;
        mem[1000] = 10'h180;
        mem[1001] = 10'h1eb;
        mem[1002] = 10'h011;
        mem[1003] = 10'h03e;
        mem[1004] = 10'h03d;
        mem[1005] = 10'h017;
        mem[1006] = 10'h000;
        mem[1007] = 10'h1d4;
        mem[1008] = 10'h00f;
        mem[1009] = 10'h08b;
        mem[1010] = 10'h37b;
        mem[1011] = 10'h0ab;
        mem[1012] = 10'h312;
        mem[1013] = 10'h373;
        mem[1014] = 10'h399;
        mem[1015] = 10'h304;
        mem[1016] = 10'h221;
        mem[1017] = 10'h39a;
        mem[1018] = 10'h3d3;
        mem[1019] = 10'h2d6;
        mem[1020] = 10'h113;
        mem[1021] = 10'h204;
        mem[1022] = 10'h055;
        mem[1023] = 10'h3a3;
    end
endmodule

module encrypt_4sbox_large8(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h3b0;
        mem[1] = 10'h205;
        mem[2] = 10'h23b;
        mem[3] = 10'h05b;
        mem[4] = 10'h0f4;
        mem[5] = 10'h398;
        mem[6] = 10'h032;
        mem[7] = 10'h002;
        mem[8] = 10'h125;
        mem[9] = 10'h2ea;
        mem[10] = 10'h280;
        mem[11] = 10'h078;
        mem[12] = 10'h3ec;
        mem[13] = 10'h2c6;
        mem[14] = 10'h124;
        mem[15] = 10'h09a;
        mem[16] = 10'h1f8;
        mem[17] = 10'h0f8;
        mem[18] = 10'h341;
        mem[19] = 10'h140;
        mem[20] = 10'h1c0;
        mem[21] = 10'h373;
        mem[22] = 10'h1d8;
        mem[23] = 10'h19a;
        mem[24] = 10'h2e9;
        mem[25] = 10'h17b;
        mem[26] = 10'h1fa;
        mem[27] = 10'h251;
        mem[28] = 10'h2ca;
        mem[29] = 10'h041;
        mem[30] = 10'h21a;
        mem[31] = 10'h03d;
        mem[32] = 10'h021;
        mem[33] = 10'h3d5;
        mem[34] = 10'h226;
        mem[35] = 10'h103;
        mem[36] = 10'h122;
        mem[37] = 10'h2b5;
        mem[38] = 10'h31f;
        mem[39] = 10'h02b;
        mem[40] = 10'h232;
        mem[41] = 10'h0ef;
        mem[42] = 10'h149;
        mem[43] = 10'h074;
        mem[44] = 10'h3bc;
        mem[45] = 10'h29e;
        mem[46] = 10'h2a9;
        mem[47] = 10'h3ce;
        mem[48] = 10'h179;
        mem[49] = 10'h0d8;
        mem[50] = 10'h220;
        mem[51] = 10'h057;
        mem[52] = 10'h119;
        mem[53] = 10'h0d9;
        mem[54] = 10'h353;
        mem[55] = 10'h120;
        mem[56] = 10'h177;
        mem[57] = 10'h1a1;
        mem[58] = 10'h176;
        mem[59] = 10'h0e9;
        mem[60] = 10'h01d;
        mem[61] = 10'h154;
        mem[62] = 10'h2b8;
        mem[63] = 10'h3bd;
        mem[64] = 10'h0d5;
        mem[65] = 10'h225;
        mem[66] = 10'h2f6;
        mem[67] = 10'h354;
        mem[68] = 10'h3ea;
        mem[69] = 10'h388;
        mem[70] = 10'h39e;
        mem[71] = 10'h2f8;
        mem[72] = 10'h11c;
        mem[73] = 10'h066;
        mem[74] = 10'h20b;
        mem[75] = 10'h247;
        mem[76] = 10'h298;
        mem[77] = 10'h18c;
        mem[78] = 10'h25e;
        mem[79] = 10'h0ee;
        mem[80] = 10'h330;
        mem[81] = 10'h051;
        mem[82] = 10'h0ba;
        mem[83] = 10'h186;
        mem[84] = 10'h3f4;
        mem[85] = 10'h234;
        mem[86] = 10'h27b;
        mem[87] = 10'h09f;
        mem[88] = 10'h067;
        mem[89] = 10'h3fd;
        mem[90] = 10'h37e;
        mem[91] = 10'h2a5;
        mem[92] = 10'h105;
        mem[93] = 10'h302;
        mem[94] = 10'h182;
        mem[95] = 10'h018;
        mem[96] = 10'h1bf;
        mem[97] = 10'h016;
        mem[98] = 10'h2f3;
        mem[99] = 10'h271;
        mem[100] = 10'h2fe;
        mem[101] = 10'h391;
        mem[102] = 10'h321;
        mem[103] = 10'h107;
        mem[104] = 10'h2b2;
        mem[105] = 10'h005;
        mem[106] = 10'h171;
        mem[107] = 10'h33a;
        mem[108] = 10'h28e;
        mem[109] = 10'h1fd;
        mem[110] = 10'h3ee;
        mem[111] = 10'h1b4;
        mem[112] = 10'h315;
        mem[113] = 10'h327;
        mem[114] = 10'h221;
        mem[115] = 10'h16b;
        mem[116] = 10'h0db;
        mem[117] = 10'h093;
        mem[118] = 10'h32c;
        mem[119] = 10'h2ef;
        mem[120] = 10'h384;
        mem[121] = 10'h030;
        mem[122] = 10'h1b1;
        mem[123] = 10'h33f;
        mem[124] = 10'h3b3;
        mem[125] = 10'h1af;
        mem[126] = 10'h29c;
        mem[127] = 10'h168;
        mem[128] = 10'h1ad;
        mem[129] = 10'h2ab;
        mem[130] = 10'h2e5;
        mem[131] = 10'h144;
        mem[132] = 10'h0bd;
        mem[133] = 10'h108;
        mem[134] = 10'h013;
        mem[135] = 10'h245;
        mem[136] = 10'h246;
        mem[137] = 10'h0bf;
        mem[138] = 10'h022;
        mem[139] = 10'h1c8;
        mem[140] = 10'h33e;
        mem[141] = 10'h0fb;
        mem[142] = 10'h101;
        mem[143] = 10'h05d;
        mem[144] = 10'h0ae;
        mem[145] = 10'h0cf;
        mem[146] = 10'h062;
        mem[147] = 10'h1cf;
        mem[148] = 10'h230;
        mem[149] = 10'h137;
        mem[150] = 10'h349;
        mem[151] = 10'h3b7;
        mem[152] = 10'h1ed;
        mem[153] = 10'h26d;
        mem[154] = 10'h02d;
        mem[155] = 10'h36b;
        mem[156] = 10'h3b4;
        mem[157] = 10'h052;
        mem[158] = 10'h39c;
        mem[159] = 10'h10c;
        mem[160] = 10'h1a3;
        mem[161] = 10'h1da;
        mem[162] = 10'h099;
        mem[163] = 10'h08e;
        mem[164] = 10'h134;
        mem[165] = 10'h023;
        mem[166] = 10'h16d;
        mem[167] = 10'h211;
        mem[168] = 10'h3b2;
        mem[169] = 10'h319;
        mem[170] = 10'h3d6;
        mem[171] = 10'h365;
        mem[172] = 10'h019;
        mem[173] = 10'h003;
        mem[174] = 10'h1b8;
        mem[175] = 10'h0a4;
        mem[176] = 10'h26c;
        mem[177] = 10'h07e;
        mem[178] = 10'h0fa;
        mem[179] = 10'h33c;
        mem[180] = 10'h340;
        mem[181] = 10'h1e0;
        mem[182] = 10'h21e;
        mem[183] = 10'h089;
        mem[184] = 10'h1f2;
        mem[185] = 10'h339;
        mem[186] = 10'h12e;
        mem[187] = 10'h377;
        mem[188] = 10'h059;
        mem[189] = 10'h0c6;
        mem[190] = 10'h025;
        mem[191] = 10'h35e;
        mem[192] = 10'h17d;
        mem[193] = 10'h2fb;
        mem[194] = 10'h3d3;
        mem[195] = 10'h0b2;
        mem[196] = 10'h20e;
        mem[197] = 10'h286;
        mem[198] = 10'h0da;
        mem[199] = 10'h32e;
        mem[200] = 10'h36f;
        mem[201] = 10'h39b;
        mem[202] = 10'h236;
        mem[203] = 10'h04b;
        mem[204] = 10'h3c6;
        mem[205] = 10'h3ed;
        mem[206] = 10'h06f;
        mem[207] = 10'h112;
        mem[208] = 10'h31e;
        mem[209] = 10'h15a;
        mem[210] = 10'h3e8;
        mem[211] = 10'h1e1;
        mem[212] = 10'h2f5;
        mem[213] = 10'h390;
        mem[214] = 10'h34d;
        mem[215] = 10'h31c;
        mem[216] = 10'h077;
        mem[217] = 10'h1a6;
        mem[218] = 10'h3e2;
        mem[219] = 10'h303;
        mem[220] = 10'h000;
        mem[221] = 10'h111;
        mem[222] = 10'h254;
        mem[223] = 10'h375;
        mem[224] = 10'h01b;
        mem[225] = 10'h2e7;
        mem[226] = 10'h2e4;
        mem[227] = 10'h329;
        mem[228] = 10'h399;
        mem[229] = 10'h212;
        mem[230] = 10'h228;
        mem[231] = 10'h1f7;
        mem[232] = 10'h1a4;
        mem[233] = 10'h100;
        mem[234] = 10'h02a;
        mem[235] = 10'h2f0;
        mem[236] = 10'h2eb;
        mem[237] = 10'h10b;
        mem[238] = 10'h3a2;
        mem[239] = 10'h300;
        mem[240] = 10'h2bb;
        mem[241] = 10'h380;
        mem[242] = 10'h033;
        mem[243] = 10'h3cc;
        mem[244] = 10'h233;
        mem[245] = 10'h02e;
        mem[246] = 10'h342;
        mem[247] = 10'h2a2;
        mem[248] = 10'h0d7;
        mem[249] = 10'h113;
        mem[250] = 10'h2ff;
        mem[251] = 10'h378;
        mem[252] = 10'h143;
        mem[253] = 10'h15b;
        mem[254] = 10'h32d;
        mem[255] = 10'h326;
        mem[256] = 10'h37c;
        mem[257] = 10'h295;
        mem[258] = 10'h22b;
        mem[259] = 10'h123;
        mem[260] = 10'h010;
        mem[261] = 10'h0b1;
        mem[262] = 10'h2ba;
        mem[263] = 10'h00d;
        mem[264] = 10'h0ce;
        mem[265] = 10'h0ed;
        mem[266] = 10'h017;
        mem[267] = 10'h381;
        mem[268] = 10'h2b7;
        mem[269] = 10'h389;
        mem[270] = 10'h0b6;
        mem[271] = 10'h364;
        mem[272] = 10'h13a;
        mem[273] = 10'h071;
        mem[274] = 10'h3fb;
        mem[275] = 10'h1ee;
        mem[276] = 10'h1f3;
        mem[277] = 10'h3bb;
        mem[278] = 10'h1d5;
        mem[279] = 10'h0d2;
        mem[280] = 10'h0ad;
        mem[281] = 10'h129;
        mem[282] = 10'h3c0;
        mem[283] = 10'h05e;
        mem[284] = 10'h3ba;
        mem[285] = 10'h310;
        mem[286] = 10'h26e;
        mem[287] = 10'h277;
        mem[288] = 10'h185;
        mem[289] = 10'h0b7;
        mem[290] = 10'h150;
        mem[291] = 10'h00f;
        mem[292] = 10'h19b;
        mem[293] = 10'h156;
        mem[294] = 10'h1fe;
        mem[295] = 10'h2d5;
        mem[296] = 10'h21d;
        mem[297] = 10'h03e;
        mem[298] = 10'h3c3;
        mem[299] = 10'h1c9;
        mem[300] = 10'h1d6;
        mem[301] = 10'h3e3;
        mem[302] = 10'h37b;
        mem[303] = 10'h044;
        mem[304] = 10'h12a;
        mem[305] = 10'h2bd;
        mem[306] = 10'h142;
        mem[307] = 10'h2fa;
        mem[308] = 10'h311;
        mem[309] = 10'h3da;
        mem[310] = 10'h12b;
        mem[311] = 10'h047;
        mem[312] = 10'h1d1;
        mem[313] = 10'h0ea;
        mem[314] = 10'h130;
        mem[315] = 10'h2d9;
        mem[316] = 10'h1a9;
        mem[317] = 10'h2cd;
        mem[318] = 10'h11f;
        mem[319] = 10'h079;
        mem[320] = 10'h133;
        mem[321] = 10'h1df;
        mem[322] = 10'h3b1;
        mem[323] = 10'h37f;
        mem[324] = 10'h0c4;
        mem[325] = 10'h1dd;
        mem[326] = 10'h2ce;
        mem[327] = 10'h36c;
        mem[328] = 10'h158;
        mem[329] = 10'h238;
        mem[330] = 10'h3a7;
        mem[331] = 10'h0a6;
        mem[332] = 10'h0a2;
        mem[333] = 10'h073;
        mem[334] = 10'h210;
        mem[335] = 10'h314;
        mem[336] = 10'h25b;
        mem[337] = 10'h2a0;
        mem[338] = 10'h00b;
        mem[339] = 10'h371;
        mem[340] = 10'h060;
        mem[341] = 10'h287;
        mem[342] = 10'h11a;
        mem[343] = 10'h114;
        mem[344] = 10'h0de;
        mem[345] = 10'h28a;
        mem[346] = 10'h191;
        mem[347] = 10'h2d7;
        mem[348] = 10'h36a;
        mem[349] = 10'h153;
        mem[350] = 10'h345;
        mem[351] = 10'h165;
        mem[352] = 10'h207;
        mem[353] = 10'h12f;
        mem[354] = 10'h1d3;
        mem[355] = 10'h020;
        mem[356] = 10'h039;
        mem[357] = 10'h0f9;
        mem[358] = 10'h3f2;
        mem[359] = 10'h0c5;
        mem[360] = 10'h28f;
        mem[361] = 10'h19c;
        mem[362] = 10'h1ec;
        mem[363] = 10'h011;
        mem[364] = 10'h370;
        mem[365] = 10'h2a3;
        mem[366] = 10'h202;
        mem[367] = 10'h23e;
        mem[368] = 10'h3e1;
        mem[369] = 10'h322;
        mem[370] = 10'h24d;
        mem[371] = 10'h087;
        mem[372] = 10'h18a;
        mem[373] = 10'h0cd;
        mem[374] = 10'h27d;
        mem[375] = 10'h1e7;
        mem[376] = 10'h35b;
        mem[377] = 10'h24a;
        mem[378] = 10'h2a6;
        mem[379] = 10'h08d;
        mem[380] = 10'h3a0;
        mem[381] = 10'h3c5;
        mem[382] = 10'h070;
        mem[383] = 10'h1e6;
        mem[384] = 10'h20a;
        mem[385] = 10'h20d;
        mem[386] = 10'h34c;
        mem[387] = 10'h0e7;
        mem[388] = 10'h34b;
        mem[389] = 10'h1b0;
        mem[390] = 10'h372;
        mem[391] = 10'h29f;
        mem[392] = 10'h324;
        mem[393] = 10'h383;
        mem[394] = 10'h009;
        mem[395] = 10'h15c;
        mem[396] = 10'h23a;
        mem[397] = 10'h2fd;
        mem[398] = 10'h260;
        mem[399] = 10'h080;
        mem[400] = 10'h1b9;
        mem[401] = 10'h1b6;
        mem[402] = 10'h17c;
        mem[403] = 10'h27a;
        mem[404] = 10'h1d9;
        mem[405] = 10'h374;
        mem[406] = 10'h14d;
        mem[407] = 10'h043;
        mem[408] = 10'h11d;
        mem[409] = 10'h36e;
        mem[410] = 10'h2d6;
        mem[411] = 10'h239;
        mem[412] = 10'h085;
        mem[413] = 10'h24b;
        mem[414] = 10'h338;
        mem[415] = 10'h036;
        mem[416] = 10'h3b8;
        mem[417] = 10'h29d;
        mem[418] = 10'h335;
        mem[419] = 10'h309;
        mem[420] = 10'h1dc;
        mem[421] = 10'h1ab;
        mem[422] = 10'h22d;
        mem[423] = 10'h046;
        mem[424] = 10'h3a4;
        mem[425] = 10'h0f7;
        mem[426] = 10'h2e8;
        mem[427] = 10'h15d;
        mem[428] = 10'h2b0;
        mem[429] = 10'h346;
        mem[430] = 10'h195;
        mem[431] = 10'h3f1;
        mem[432] = 10'h2d8;
        mem[433] = 10'h386;
        mem[434] = 10'h3e4;
        mem[435] = 10'h07a;
        mem[436] = 10'h356;
        mem[437] = 10'h3ad;
        mem[438] = 10'h3fa;
        mem[439] = 10'h235;
        mem[440] = 10'h36d;
        mem[441] = 10'h068;
        mem[442] = 10'h2cf;
        mem[443] = 10'h25f;
        mem[444] = 10'h3c4;
        mem[445] = 10'h0ff;
        mem[446] = 10'h2af;
        mem[447] = 10'h082;
        mem[448] = 10'h268;
        mem[449] = 10'h242;
        mem[450] = 10'h2b9;
        mem[451] = 10'h332;
        mem[452] = 10'h2c8;
        mem[453] = 10'h2b1;
        mem[454] = 10'h28b;
        mem[455] = 10'h252;
        mem[456] = 10'h334;
        mem[457] = 10'h3c8;
        mem[458] = 10'h2ec;
        mem[459] = 10'h259;
        mem[460] = 10'h164;
        mem[461] = 10'h214;
        mem[462] = 10'h04f;
        mem[463] = 10'h253;
        mem[464] = 10'h3c7;
        mem[465] = 10'h07d;
        mem[466] = 10'h0f3;
        mem[467] = 10'h284;
        mem[468] = 10'h1e2;
        mem[469] = 10'h135;
        mem[470] = 10'h0b9;
        mem[471] = 10'h0a1;
        mem[472] = 10'h33d;
        mem[473] = 10'h050;
        mem[474] = 10'h1c2;
        mem[475] = 10'h2e6;
        mem[476] = 10'h15e;
        mem[477] = 10'h394;
        mem[478] = 10'h083;
        mem[479] = 10'h159;
        mem[480] = 10'h00e;
        mem[481] = 10'h13d;
        mem[482] = 10'h03f;
        mem[483] = 10'h1f9;
        mem[484] = 10'h2d0;
        mem[485] = 10'h172;
        mem[486] = 10'h2c7;
        mem[487] = 10'h2f4;
        mem[488] = 10'h05a;
        mem[489] = 10'h21b;
        mem[490] = 10'h2f7;
        mem[491] = 10'h2c0;
        mem[492] = 10'h16c;
        mem[493] = 10'h24c;
        mem[494] = 10'h3e5;
        mem[495] = 10'h086;
        mem[496] = 10'h2cc;
        mem[497] = 10'h38a;
        mem[498] = 10'h273;
        mem[499] = 10'h320;
        mem[500] = 10'h209;
        mem[501] = 10'h0a3;
        mem[502] = 10'h358;
        mem[503] = 10'h2c3;
        mem[504] = 10'h1a8;
        mem[505] = 10'h037;
        mem[506] = 10'h027;
        mem[507] = 10'h0d1;
        mem[508] = 10'h38e;
        mem[509] = 10'h387;
        mem[510] = 10'h163;
        mem[511] = 10'h25c;
        mem[512] = 10'h3d0;
        mem[513] = 10'h313;
        mem[514] = 10'h1cd;
        mem[515] = 10'h10e;
        mem[516] = 10'h199;
        mem[517] = 10'h30b;
        mem[518] = 10'h06a;
        mem[519] = 10'h0df;
        mem[520] = 10'h2a1;
        mem[521] = 10'h3d4;
        mem[522] = 10'h282;
        mem[523] = 10'h3fe;
        mem[524] = 10'h06b;
        mem[525] = 10'h2c9;
        mem[526] = 10'h337;
        mem[527] = 10'h2d2;
        mem[528] = 10'h31a;
        mem[529] = 10'h094;
        mem[530] = 10'h0e1;
        mem[531] = 10'h075;
        mem[532] = 10'h007;
        mem[533] = 10'h01a;
        mem[534] = 10'h0ab;
        mem[535] = 10'h004;
        mem[536] = 10'h2bf;
        mem[537] = 10'h19e;
        mem[538] = 10'h29a;
        mem[539] = 10'h126;
        mem[540] = 10'h141;
        mem[541] = 10'h116;
        mem[542] = 10'h1cb;
        mem[543] = 10'h362;
        mem[544] = 10'h1d7;
        mem[545] = 10'h396;
        mem[546] = 10'h06e;
        mem[547] = 10'h283;
        mem[548] = 10'h2b3;
        mem[549] = 10'h3eb;
        mem[550] = 10'h222;
        mem[551] = 10'h1e3;
        mem[552] = 10'h376;
        mem[553] = 10'h34e;
        mem[554] = 10'h312;
        mem[555] = 10'h3ef;
        mem[556] = 10'h2f9;
        mem[557] = 10'h1a7;
        mem[558] = 10'h1e5;
        mem[559] = 10'h0f6;
        mem[560] = 10'h157;
        mem[561] = 10'h187;
        mem[562] = 10'h18e;
        mem[563] = 10'h155;
        mem[564] = 10'h30a;
        mem[565] = 10'h363;
        mem[566] = 10'h265;
        mem[567] = 10'h0dc;
        mem[568] = 10'h1a2;
        mem[569] = 10'h3c2;
        mem[570] = 10'h1b3;
        mem[571] = 10'h3b9;
        mem[572] = 10'h2e3;
        mem[573] = 10'h2ee;
        mem[574] = 10'h1cc;
        mem[575] = 10'h19d;
        mem[576] = 10'h270;
        mem[577] = 10'h145;
        mem[578] = 10'h258;
        mem[579] = 10'h229;
        mem[580] = 10'h227;
        mem[581] = 10'h2db;
        mem[582] = 10'h131;
        mem[583] = 10'h04e;
        mem[584] = 10'h333;
        mem[585] = 10'h1fc;
        mem[586] = 10'h1e4;
        mem[587] = 10'h05f;
        mem[588] = 10'h359;
        mem[589] = 10'h2d1;
        mem[590] = 10'h216;
        mem[591] = 10'h276;
        mem[592] = 10'h24f;
        mem[593] = 10'h0e3;
        mem[594] = 10'h2d4;
        mem[595] = 10'h3a5;
        mem[596] = 10'h098;
        mem[597] = 10'h325;
        mem[598] = 10'h3e7;
        mem[599] = 10'h301;
        mem[600] = 10'h3cf;
        mem[601] = 10'h181;
        mem[602] = 10'h344;
        mem[603] = 10'h2c2;
        mem[604] = 10'h317;
        mem[605] = 10'h30c;
        mem[606] = 10'h290;
        mem[607] = 10'h024;
        mem[608] = 10'h096;
        mem[609] = 10'h316;
        mem[610] = 10'h2bc;
        mem[611] = 10'h3ae;
        mem[612] = 10'h1c5;
        mem[613] = 10'h2de;
        mem[614] = 10'h30e;
        mem[615] = 10'h2fc;
        mem[616] = 10'h03a;
        mem[617] = 10'h1ff;
        mem[618] = 10'h13e;
        mem[619] = 10'h29b;
        mem[620] = 10'h3dc;
        mem[621] = 10'h1f1;
        mem[622] = 10'h30d;
        mem[623] = 10'h1db;
        mem[624] = 10'h257;
        mem[625] = 10'h063;
        mem[626] = 10'h21f;
        mem[627] = 10'h1c7;
        mem[628] = 10'h2a4;
        mem[629] = 10'h256;
        mem[630] = 10'h351;
        mem[631] = 10'h1e8;
        mem[632] = 10'h01c;
        mem[633] = 10'h034;
        mem[634] = 10'h048;
        mem[635] = 10'h35a;
        mem[636] = 10'h128;
        mem[637] = 10'h0e4;
        mem[638] = 10'h32f;
        mem[639] = 10'h147;
        mem[640] = 10'h291;
        mem[641] = 10'h1c6;
        mem[642] = 10'h072;
        mem[643] = 10'h2b6;
        mem[644] = 10'h3f9;
        mem[645] = 10'h097;
        mem[646] = 10'h22f;
        mem[647] = 10'h244;
        mem[648] = 10'h1be;
        mem[649] = 10'h194;
        mem[650] = 10'h0eb;
        mem[651] = 10'h1bd;
        mem[652] = 10'h188;
        mem[653] = 10'h091;
        mem[654] = 10'h0e2;
        mem[655] = 10'h3ab;
        mem[656] = 10'h102;
        mem[657] = 10'h33b;
        mem[658] = 10'h139;
        mem[659] = 10'h38b;
        mem[660] = 10'h1de;
        mem[661] = 10'h10a;
        mem[662] = 10'h042;
        mem[663] = 10'h203;
        mem[664] = 10'h1bc;
        mem[665] = 10'h343;
        mem[666] = 10'h061;
        mem[667] = 10'h008;
        mem[668] = 10'h1a0;
        mem[669] = 10'h26f;
        mem[670] = 10'h0b0;
        mem[671] = 10'h304;
        mem[672] = 10'h084;
        mem[673] = 10'h045;
        mem[674] = 10'h223;
        mem[675] = 10'h279;
        mem[676] = 10'h192;
        mem[677] = 10'h248;
        mem[678] = 10'h1b2;
        mem[679] = 10'h224;
        mem[680] = 10'h2f2;
        mem[681] = 10'h169;
        mem[682] = 10'h3df;
        mem[683] = 10'h266;
        mem[684] = 10'h272;
        mem[685] = 10'h281;
        mem[686] = 10'h1d2;
        mem[687] = 10'h146;
        mem[688] = 10'h088;
        mem[689] = 10'h3fc;
        mem[690] = 10'h028;
        mem[691] = 10'h0f5;
        mem[692] = 10'h2df;
        mem[693] = 10'h385;
        mem[694] = 10'h160;
        mem[695] = 10'h255;
        mem[696] = 10'h07b;
        mem[697] = 10'h293;
        mem[698] = 10'h3e6;
        mem[699] = 10'h3f8;
        mem[700] = 10'h184;
        mem[701] = 10'h1d4;
        mem[702] = 10'h180;
        mem[703] = 10'h2cb;
        mem[704] = 10'h3b6;
        mem[705] = 10'h1c3;
        mem[706] = 10'h0c9;
        mem[707] = 10'h17a;
        mem[708] = 10'h393;
        mem[709] = 10'h069;
        mem[710] = 10'h0b8;
        mem[711] = 10'h3a3;
        mem[712] = 10'h189;
        mem[713] = 10'h0a9;
        mem[714] = 10'h37a;
        mem[715] = 10'h1ef;
        mem[716] = 10'h0c7;
        mem[717] = 10'h0fd;
        mem[718] = 10'h0af;
        mem[719] = 10'h198;
        mem[720] = 10'h18f;
        mem[721] = 10'h264;
        mem[722] = 10'h13b;
        mem[723] = 10'h136;
        mem[724] = 10'h06c;
        mem[725] = 10'h269;
        mem[726] = 10'h215;
        mem[727] = 10'h0a8;
        mem[728] = 10'h288;
        mem[729] = 10'h06d;
        mem[730] = 10'h336;
        mem[731] = 10'h03b;
        mem[732] = 10'h0e5;
        mem[733] = 10'h081;
        mem[734] = 10'h3a6;
        mem[735] = 10'h0a0;
        mem[736] = 10'h08c;
        mem[737] = 10'h237;
        mem[738] = 10'h190;
        mem[739] = 10'h1b7;
        mem[740] = 10'h243;
        mem[741] = 10'h3af;
        mem[742] = 10'h0aa;
        mem[743] = 10'h3a9;
        mem[744] = 10'h38d;
        mem[745] = 10'h01e;
        mem[746] = 10'h055;
        mem[747] = 10'h173;
        mem[748] = 10'h348;
        mem[749] = 10'h22a;
        mem[750] = 10'h1c4;
        mem[751] = 10'h058;
        mem[752] = 10'h2be;
        mem[753] = 10'h0bb;
        mem[754] = 10'h0bc;
        mem[755] = 10'h0fc;
        mem[756] = 10'h1e9;
        mem[757] = 10'h0ec;
        mem[758] = 10'h0f0;
        mem[759] = 10'h3bf;
        mem[760] = 10'h121;
        mem[761] = 10'h3c9;
        mem[762] = 10'h04a;
        mem[763] = 10'h26a;
        mem[764] = 10'h11e;
        mem[765] = 10'h09e;
        mem[766] = 10'h3be;
        mem[767] = 10'h367;
        mem[768] = 10'h2da;
        mem[769] = 10'h28c;
        mem[770] = 10'h0c2;
        mem[771] = 10'h379;
        mem[772] = 10'h1aa;
        mem[773] = 10'h397;
        mem[774] = 10'h0c3;
        mem[775] = 10'h31b;
        mem[776] = 10'h2ac;
        mem[777] = 10'h092;
        mem[778] = 10'h0fe;
        mem[779] = 10'h152;
        mem[780] = 10'h0b3;
        mem[781] = 10'h0d0;
        mem[782] = 10'h1d0;
        mem[783] = 10'h217;
        mem[784] = 10'h328;
        mem[785] = 10'h240;
        mem[786] = 10'h16f;
        mem[787] = 10'h1ba;
        mem[788] = 10'h1f0;
        mem[789] = 10'h323;
        mem[790] = 10'h09c;
        mem[791] = 10'h2dd;
        mem[792] = 10'h095;
        mem[793] = 10'h2e2;
        mem[794] = 10'h109;
        mem[795] = 10'h1ea;
        mem[796] = 10'h25a;
        mem[797] = 10'h14b;
        mem[798] = 10'h015;
        mem[799] = 10'h1ca;
        mem[800] = 10'h006;
        mem[801] = 10'h2c5;
        mem[802] = 10'h183;
        mem[803] = 10'h307;
        mem[804] = 10'h0ac;
        mem[805] = 10'h22c;
        mem[806] = 10'h3d2;
        mem[807] = 10'h10d;
        mem[808] = 10'h30f;
        mem[809] = 10'h285;
        mem[810] = 10'h2dc;
        mem[811] = 10'h2b4;
        mem[812] = 10'h0dd;
        mem[813] = 10'h076;
        mem[814] = 10'h00c;
        mem[815] = 10'h2aa;
        mem[816] = 10'h174;
        mem[817] = 10'h3f6;
        mem[818] = 10'h263;
        mem[819] = 10'h090;
        mem[820] = 10'h11b;
        mem[821] = 10'h110;
        mem[822] = 10'h241;
        mem[823] = 10'h249;
        mem[824] = 10'h104;
        mem[825] = 10'h294;
        mem[826] = 10'h275;
        mem[827] = 10'h204;
        mem[828] = 10'h106;
        mem[829] = 10'h35c;
        mem[830] = 10'h331;
        mem[831] = 10'h20f;
        mem[832] = 10'h2c1;
        mem[833] = 10'h3de;
        mem[834] = 10'h01f;
        mem[835] = 10'h08b;
        mem[836] = 10'h274;
        mem[837] = 10'h262;
        mem[838] = 10'h382;
        mem[839] = 10'h132;
        mem[840] = 10'h37d;
        mem[841] = 10'h267;
        mem[842] = 10'h10f;
        mem[843] = 10'h218;
        mem[844] = 10'h0a7;
        mem[845] = 10'h3ff;
        mem[846] = 10'h0c8;
        mem[847] = 10'h1f4;
        mem[848] = 10'h040;
        mem[849] = 10'h2e1;
        mem[850] = 10'h05c;
        mem[851] = 10'h15f;
        mem[852] = 10'h231;
        mem[853] = 10'h289;
        mem[854] = 10'h14f;
        mem[855] = 10'h17f;
        mem[856] = 10'h2a7;
        mem[857] = 10'h3d1;
        mem[858] = 10'h392;
        mem[859] = 10'h18b;
        mem[860] = 10'h3dd;
        mem[861] = 10'h3f7;
        mem[862] = 10'h34f;
        mem[863] = 10'h3f5;
        mem[864] = 10'h16a;
        mem[865] = 10'h299;
        mem[866] = 10'h278;
        mem[867] = 10'h0be;
        mem[868] = 10'h3e0;
        mem[869] = 10'h08a;
        mem[870] = 10'h38c;
        mem[871] = 10'h035;
        mem[872] = 10'h04d;
        mem[873] = 10'h3cd;
        mem[874] = 10'h064;
        mem[875] = 10'h029;
        mem[876] = 10'h308;
        mem[877] = 10'h1f6;
        mem[878] = 10'h07c;
        mem[879] = 10'h16e;
        mem[880] = 10'h39f;
        mem[881] = 10'h3ac;
        mem[882] = 10'h0a5;
        mem[883] = 10'h14e;
        mem[884] = 10'h305;
        mem[885] = 10'h368;
        mem[886] = 10'h3e9;
        mem[887] = 10'h193;
        mem[888] = 10'h09d;
        mem[889] = 10'h23f;
        mem[890] = 10'h3a1;
        mem[891] = 10'h3f0;
        mem[892] = 10'h197;
        mem[893] = 10'h0c0;
        mem[894] = 10'h200;
        mem[895] = 10'h361;
        mem[896] = 10'h08f;
        mem[897] = 10'h053;
        mem[898] = 10'h0ca;
        mem[899] = 10'h3c1;
        mem[900] = 10'h3b5;
        mem[901] = 10'h161;
        mem[902] = 10'h038;
        mem[903] = 10'h166;
        mem[904] = 10'h3d9;
        mem[905] = 10'h178;
        mem[906] = 10'h02c;
        mem[907] = 10'h18d;
        mem[908] = 10'h201;
        mem[909] = 10'h031;
        mem[910] = 10'h2f1;
        mem[911] = 10'h28d;
        mem[912] = 10'h127;
        mem[913] = 10'h1f5;
        mem[914] = 10'h3db;
        mem[915] = 10'h20c;
        mem[916] = 10'h25d;
        mem[917] = 10'h2e0;
        mem[918] = 10'h02f;
        mem[919] = 10'h2ae;
        mem[920] = 10'h395;
        mem[921] = 10'h1ae;
        mem[922] = 10'h219;
        mem[923] = 10'h00a;
        mem[924] = 10'h170;
        mem[925] = 10'h0d4;
        mem[926] = 10'h0e0;
        mem[927] = 10'h117;
        mem[928] = 10'h148;
        mem[929] = 10'h17e;
        mem[930] = 10'h162;
        mem[931] = 10'h350;
        mem[932] = 10'h1b5;
        mem[933] = 10'h32b;
        mem[934] = 10'h0f1;
        mem[935] = 10'h012;
        mem[936] = 10'h35d;
        mem[937] = 10'h31d;
        mem[938] = 10'h151;
        mem[939] = 10'h26b;
        mem[940] = 10'h0d6;
        mem[941] = 10'h2a8;
        mem[942] = 10'h014;
        mem[943] = 10'h38f;
        mem[944] = 10'h2d3;
        mem[945] = 10'h12c;
        mem[946] = 10'h366;
        mem[947] = 10'h056;
        mem[948] = 10'h3aa;
        mem[949] = 10'h1ac;
        mem[950] = 10'h292;
        mem[951] = 10'h2c4;
        mem[952] = 10'h3f3;
        mem[953] = 10'h0d3;
        mem[954] = 10'h213;
        mem[955] = 10'h22e;
        mem[956] = 10'h049;
        mem[957] = 10'h03c;
        mem[958] = 10'h35f;
        mem[959] = 10'h13f;
        mem[960] = 10'h39d;
        mem[961] = 10'h24e;
        mem[962] = 10'h1fb;
        mem[963] = 10'h0c1;
        mem[964] = 10'h115;
        mem[965] = 10'h1bb;
        mem[966] = 10'h2ed;
        mem[967] = 10'h04c;
        mem[968] = 10'h27e;
        mem[969] = 10'h250;
        mem[970] = 10'h001;
        mem[971] = 10'h318;
        mem[972] = 10'h1eb;
        mem[973] = 10'h357;
        mem[974] = 10'h167;
        mem[975] = 10'h347;
        mem[976] = 10'h19f;
        mem[977] = 10'h026;
        mem[978] = 10'h297;
        mem[979] = 10'h2ad;
        mem[980] = 10'h39a;
        mem[981] = 10'h3ca;
        mem[982] = 10'h352;
        mem[983] = 10'h196;
        mem[984] = 10'h261;
        mem[985] = 10'h3d7;
        mem[986] = 10'h1c1;
        mem[987] = 10'h138;
        mem[988] = 10'h14c;
        mem[989] = 10'h13c;
        mem[990] = 10'h21c;
        mem[991] = 10'h369;
        mem[992] = 10'h23c;
        mem[993] = 10'h360;
        mem[994] = 10'h355;
        mem[995] = 10'h175;
        mem[996] = 10'h0cb;
        mem[997] = 10'h27c;
        mem[998] = 10'h34a;
        mem[999] = 10'h1ce;
        mem[1000] = 10'h118;
        mem[1001] = 10'h0e6;
        mem[1002] = 10'h3d8;
        mem[1003] = 10'h0f2;
        mem[1004] = 10'h09b;
        mem[1005] = 10'h27f;
        mem[1006] = 10'h12d;
        mem[1007] = 10'h1a5;
        mem[1008] = 10'h0e8;
        mem[1009] = 10'h3cb;
        mem[1010] = 10'h0b5;
        mem[1011] = 10'h065;
        mem[1012] = 10'h206;
        mem[1013] = 10'h0cc;
        mem[1014] = 10'h14a;
        mem[1015] = 10'h306;
        mem[1016] = 10'h0b4;
        mem[1017] = 10'h23d;
        mem[1018] = 10'h07f;
        mem[1019] = 10'h054;
        mem[1020] = 10'h296;
        mem[1021] = 10'h32a;
        mem[1022] = 10'h208;
        mem[1023] = 10'h3a8;
    end
endmodule

module encrypt_4sbox_large9(clk, a_in, b_in, a_out, b_out);
    input clk;
    input [9:0] a_in;
    output reg [9:0] a_out;
    input [9:0] b_in;
    output reg [9:0] b_out;
    reg [9:0] mem[0:1023];
    always @(posedge clk) begin
        a_out <= mem[a_in];
        b_out <= mem[b_in];
    end
    initial begin
        mem[0] = 10'h384;
        mem[1] = 10'h328;
        mem[2] = 10'h306;
        mem[3] = 10'h05b;
        mem[4] = 10'h0de;
        mem[5] = 10'h0d2;
        mem[6] = 10'h1ce;
        mem[7] = 10'h04c;
        mem[8] = 10'h3d9;
        mem[9] = 10'h3b0;
        mem[10] = 10'h157;
        mem[11] = 10'h307;
        mem[12] = 10'h268;
        mem[13] = 10'h382;
        mem[14] = 10'h149;
        mem[15] = 10'h1ae;
        mem[16] = 10'h176;
        mem[17] = 10'h22a;
        mem[18] = 10'h03a;
        mem[19] = 10'h2b6;
        mem[20] = 10'h10c;
        mem[21] = 10'h13a;
        mem[22] = 10'h0ee;
        mem[23] = 10'h291;
        mem[24] = 10'h3c1;
        mem[25] = 10'h2ba;
        mem[26] = 10'h016;
        mem[27] = 10'h059;
        mem[28] = 10'h11f;
        mem[29] = 10'h321;
        mem[30] = 10'h0a7;
        mem[31] = 10'h2fe;
        mem[32] = 10'h287;
        mem[33] = 10'h162;
        mem[34] = 10'h35f;
        mem[35] = 10'h112;
        mem[36] = 10'h14f;
        mem[37] = 10'h350;
        mem[38] = 10'h0ff;
        mem[39] = 10'h334;
        mem[40] = 10'h141;
        mem[41] = 10'h044;
        mem[42] = 10'h058;
        mem[43] = 10'h117;
        mem[44] = 10'h3a5;
        mem[45] = 10'h045;
        mem[46] = 10'h030;
        mem[47] = 10'h2a0;
        mem[48] = 10'h2f5;
        mem[49] = 10'h39c;
        mem[50] = 10'h305;
        mem[51] = 10'h3e8;
        mem[52] = 10'h25e;
        mem[53] = 10'h2cf;
        mem[54] = 10'h3a4;
        mem[55] = 10'h368;
        mem[56] = 10'h0c6;
        mem[57] = 10'h167;
        mem[58] = 10'h3a9;
        mem[59] = 10'h0a4;
        mem[60] = 10'h0f4;
        mem[61] = 10'h271;
        mem[62] = 10'h0e1;
        mem[63] = 10'h2ac;
        mem[64] = 10'h165;
        mem[65] = 10'h163;
        mem[66] = 10'h18d;
        mem[67] = 10'h042;
        mem[68] = 10'h370;
        mem[69] = 10'h183;
        mem[70] = 10'h002;
        mem[71] = 10'h107;
        mem[72] = 10'h360;
        mem[73] = 10'h234;
        mem[74] = 10'h286;
        mem[75] = 10'h229;
        mem[76] = 10'h0ae;
        mem[77] = 10'h001;
        mem[78] = 10'h22b;
        mem[79] = 10'h2e8;
        mem[80] = 10'h30c;
        mem[81] = 10'h2e0;
        mem[82] = 10'h115;
        mem[83] = 10'h1e6;
        mem[84] = 10'h330;
        mem[85] = 10'h261;
        mem[86] = 10'h26d;
        mem[87] = 10'h2d3;
        mem[88] = 10'h26f;
        mem[89] = 10'h2b5;
        mem[90] = 10'h319;
        mem[91] = 10'h2bf;
        mem[92] = 10'h1c6;
        mem[93] = 10'h29c;
        mem[94] = 10'h1dc;
        mem[95] = 10'h237;
        mem[96] = 10'h2df;
        mem[97] = 10'h097;
        mem[98] = 10'h1a1;
        mem[99] = 10'h31f;
        mem[100] = 10'h031;
        mem[101] = 10'h2cb;
        mem[102] = 10'h053;
        mem[103] = 10'h193;
        mem[104] = 10'h03b;
        mem[105] = 10'h278;
        mem[106] = 10'h120;
        mem[107] = 10'h32d;
        mem[108] = 10'h1f5;
        mem[109] = 10'h23e;
        mem[110] = 10'h21d;
        mem[111] = 10'h200;
        mem[112] = 10'h378;
        mem[113] = 10'h0ce;
        mem[114] = 10'h3e0;
        mem[115] = 10'h0c9;
        mem[116] = 10'h0c8;
        mem[117] = 10'h0d8;
        mem[118] = 10'h14d;
        mem[119] = 10'h2c6;
        mem[120] = 10'h1f6;
        mem[121] = 10'h348;
        mem[122] = 10'h265;
        mem[123] = 10'h398;
        mem[124] = 10'h340;
        mem[125] = 10'h29f;
        mem[126] = 10'h31d;
        mem[127] = 10'h0d4;
        mem[128] = 10'h020;
        mem[129] = 10'h351;
        mem[130] = 10'h07b;
        mem[131] = 10'h01f;
        mem[132] = 10'h0f2;
        mem[133] = 10'h0a2;
        mem[134] = 10'h0e6;
        mem[135] = 10'h221;
        mem[136] = 10'h122;
        mem[137] = 10'h20e;
        mem[138] = 10'h230;
        mem[139] = 10'h263;
        mem[140] = 10'h07e;
        mem[141] = 10'h1d7;
        mem[142] = 10'h02c;
        mem[143] = 10'h2d0;
        mem[144] = 10'h3b1;
        mem[145] = 10'h0d1;
        mem[146] = 10'h15c;
        mem[147] = 10'h13b;
        mem[148] = 10'h36e;
        mem[149] = 10'h25a;
        mem[150] = 10'h39f;
        mem[151] = 10'h214;
        mem[152] = 10'h31a;
        mem[153] = 10'h1ab;
        mem[154] = 10'h353;
        mem[155] = 10'h07f;
        mem[156] = 10'h2dd;
        mem[157] = 10'h12b;
        mem[158] = 10'h217;
        mem[159] = 10'h223;
        mem[160] = 10'h32a;
        mem[161] = 10'h04d;
        mem[162] = 10'h20c;
        mem[163] = 10'h20f;
        mem[164] = 10'h049;
        mem[165] = 10'h0d0;
        mem[166] = 10'h178;
        mem[167] = 10'h139;
        mem[168] = 10'h2f0;
        mem[169] = 10'h20d;
        mem[170] = 10'h02f;
        mem[171] = 10'h272;
        mem[172] = 10'h3e5;
        mem[173] = 10'h025;
        mem[174] = 10'h2d7;
        mem[175] = 10'h2c9;
        mem[176] = 10'h23a;
        mem[177] = 10'h088;
        mem[178] = 10'h1fe;
        mem[179] = 10'h155;
        mem[180] = 10'h147;
        mem[181] = 10'h156;
        mem[182] = 10'h0a9;
        mem[183] = 10'h253;
        mem[184] = 10'h3b9;
        mem[185] = 10'h1ec;
        mem[186] = 10'h1d3;
        mem[187] = 10'h366;
        mem[188] = 10'h339;
        mem[189] = 10'h3ad;
        mem[190] = 10'h177;
        mem[191] = 10'h0f0;
        mem[192] = 10'h3cd;
        mem[193] = 10'h346;
        mem[194] = 10'h35d;
        mem[195] = 10'h17d;
        mem[196] = 10'h085;
        mem[197] = 10'h3c2;
        mem[198] = 10'h05d;
        mem[199] = 10'h26a;
        mem[200] = 10'h3f0;
        mem[201] = 10'h326;
        mem[202] = 10'h28d;
        mem[203] = 10'h0da;
        mem[204] = 10'h021;
        mem[205] = 10'h173;
        mem[206] = 10'h161;
        mem[207] = 10'h2ed;
        mem[208] = 10'h15d;
        mem[209] = 10'h094;
        mem[210] = 10'h0a1;
        mem[211] = 10'h1ad;
        mem[212] = 10'h074;
        mem[213] = 10'h2ab;
        mem[214] = 10'h196;
        mem[215] = 10'h37a;
        mem[216] = 10'h061;
        mem[217] = 10'h06a;
        mem[218] = 10'h1d9;
        mem[219] = 10'h014;
        mem[220] = 10'h17c;
        mem[221] = 10'h103;
        mem[222] = 10'h38c;
        mem[223] = 10'h1b4;
        mem[224] = 10'h30f;
        mem[225] = 10'h136;
        mem[226] = 10'h209;
        mem[227] = 10'h2ff;
        mem[228] = 10'h31c;
        mem[229] = 10'h3c9;
        mem[230] = 10'h0f5;
        mem[231] = 10'h332;
        mem[232] = 10'h1a8;
        mem[233] = 10'h2bd;
        mem[234] = 10'h345;
        mem[235] = 10'h0bc;
        mem[236] = 10'h089;
        mem[237] = 10'h29d;
        mem[238] = 10'h073;
        mem[239] = 10'h39b;
        mem[240] = 10'h0cb;
        mem[241] = 10'h34f;
        mem[242] = 10'h038;
        mem[243] = 10'h2ec;
        mem[244] = 10'h154;
        mem[245] = 10'h241;
        mem[246] = 10'h201;
        mem[247] = 10'h1fc;
        mem[248] = 10'h2a2;
        mem[249] = 10'h28a;
        mem[250] = 10'h015;
        mem[251] = 10'h1c0;
        mem[252] = 10'h1d0;
        mem[253] = 10'h37b;
        mem[254] = 10'h248;
        mem[255] = 10'h1e7;
        mem[256] = 10'h080;
        mem[257] = 10'h2cd;
        mem[258] = 10'h239;
        mem[259] = 10'h33d;
        mem[260] = 10'h1d6;
        mem[261] = 10'h298;
        mem[262] = 10'h06f;
        mem[263] = 10'h30e;
        mem[264] = 10'h1ba;
        mem[265] = 10'h1f1;
        mem[266] = 10'h064;
        mem[267] = 10'h078;
        mem[268] = 10'h39e;
        mem[269] = 10'h3ee;
        mem[270] = 10'h187;
        mem[271] = 10'h3c8;
        mem[272] = 10'h212;
        mem[273] = 10'h1b9;
        mem[274] = 10'h2b3;
        mem[275] = 10'h3aa;
        mem[276] = 10'h3f8;
        mem[277] = 10'h1b0;
        mem[278] = 10'h39d;
        mem[279] = 10'h2eb;
        mem[280] = 10'h205;
        mem[281] = 10'h04a;
        mem[282] = 10'h260;
        mem[283] = 10'h0bd;
        mem[284] = 10'h381;
        mem[285] = 10'h086;
        mem[286] = 10'h3e1;
        mem[287] = 10'h3ec;
        mem[288] = 10'h2dc;
        mem[289] = 10'h2a4;
        mem[290] = 10'h22c;
        mem[291] = 10'h22d;
        mem[292] = 10'h2e7;
        mem[293] = 10'h0fc;
        mem[294] = 10'h374;
        mem[295] = 10'h179;
        mem[296] = 10'h124;
        mem[297] = 10'h0b0;
        mem[298] = 10'h1d4;
        mem[299] = 10'h28e;
        mem[300] = 10'h1e2;
        mem[301] = 10'h2b0;
        mem[302] = 10'h3fd;
        mem[303] = 10'h3ba;
        mem[304] = 10'h376;
        mem[305] = 10'h0af;
        mem[306] = 10'h03f;
        mem[307] = 10'h30b;
        mem[308] = 10'h18c;
        mem[309] = 10'h232;
        mem[310] = 10'h130;
        mem[311] = 10'h3e6;
        mem[312] = 10'h2f4;
        mem[313] = 10'h1ee;
        mem[314] = 10'h0c7;
        mem[315] = 10'h151;
        mem[316] = 10'h28f;
        mem[317] = 10'h056;
        mem[318] = 10'h1dd;
        mem[319] = 10'h2f2;
        mem[320] = 10'h14e;
        mem[321] = 10'h20a;
        mem[322] = 10'h2b9;
        mem[323] = 10'h2e3;
        mem[324] = 10'h134;
        mem[325] = 10'h3d1;
        mem[326] = 10'h27e;
        mem[327] = 10'h0c2;
        mem[328] = 10'h005;
        mem[329] = 10'h1a0;
        mem[330] = 10'h3f7;
        mem[331] = 10'h1c5;
        mem[332] = 10'h3b7;
        mem[333] = 10'h3cc;
        mem[334] = 10'h24d;
        mem[335] = 10'h03c;
        mem[336] = 10'h19a;
        mem[337] = 10'h023;
        mem[338] = 10'h343;
        mem[339] = 10'h076;
        mem[340] = 10'h1d8;
        mem[341] = 10'h3b6;
        mem[342] = 10'h0b8;
        mem[343] = 10'h36d;
        mem[344] = 10'h392;
        mem[345] = 10'h1a4;
        mem[346] = 10'h040;
        mem[347] = 10'h17f;
        mem[348] = 10'h121;
        mem[349] = 10'h2ae;
        mem[350] = 10'h132;
        mem[351] = 10'h397;
        mem[352] = 10'h11e;
        mem[353] = 10'h37e;
        mem[354] = 10'h1ac;
        mem[355] = 10'h222;
        mem[356] = 10'h3c4;
        mem[357] = 10'h1bc;
        mem[358] = 10'h123;
        mem[359] = 10'h2c2;
        mem[360] = 10'h08d;
        mem[361] = 10'h0b1;
        mem[362] = 10'h341;
        mem[363] = 10'h1a2;
        mem[364] = 10'h258;
        mem[365] = 10'h164;
        mem[366] = 10'h12c;
        mem[367] = 10'h0b7;
        mem[368] = 10'h3ab;
        mem[369] = 10'h363;
        mem[370] = 10'h2e5;
        mem[371] = 10'h09f;
        mem[372] = 10'h0dd;
        mem[373] = 10'h0a8;
        mem[374] = 10'h1d1;
        mem[375] = 10'h2f8;
        mem[376] = 10'h104;
        mem[377] = 10'h2e9;
        mem[378] = 10'h22e;
        mem[379] = 10'h3f4;
        mem[380] = 10'h0e3;
        mem[381] = 10'h116;
        mem[382] = 10'h27f;
        mem[383] = 10'h102;
        mem[384] = 10'h304;
        mem[385] = 10'h13c;
        mem[386] = 10'h1ef;
        mem[387] = 10'h08b;
        mem[388] = 10'h293;
        mem[389] = 10'h2f7;
        mem[390] = 10'h228;
        mem[391] = 10'h06d;
        mem[392] = 10'h365;
        mem[393] = 10'h309;
        mem[394] = 10'h349;
        mem[395] = 10'h2f3;
        mem[396] = 10'h00a;
        mem[397] = 10'h240;
        mem[398] = 10'h18f;
        mem[399] = 10'h20b;
        mem[400] = 10'h1e8;
        mem[401] = 10'h05e;
        mem[402] = 10'h3f1;
        mem[403] = 10'h138;
        mem[404] = 10'h093;
        mem[405] = 10'h11d;
        mem[406] = 10'h135;
        mem[407] = 10'h259;
        mem[408] = 10'h210;
        mem[409] = 10'h3da;
        mem[410] = 10'h0c4;
        mem[411] = 10'h213;
        mem[412] = 10'h043;
        mem[413] = 10'h0b6;
        mem[414] = 10'h2fd;
        mem[415] = 10'h19f;
        mem[416] = 10'h2c1;
        mem[417] = 10'h000;
        mem[418] = 10'h2a7;
        mem[419] = 10'h3a7;
        mem[420] = 10'h0a3;
        mem[421] = 10'h3be;
        mem[422] = 10'h2c3;
        mem[423] = 10'h10b;
        mem[424] = 10'h2a6;
        mem[425] = 10'h096;
        mem[426] = 10'h0d3;
        mem[427] = 10'h275;
        mem[428] = 10'h3a3;
        mem[429] = 10'h359;
        mem[430] = 10'h358;
        mem[431] = 10'h1f8;
        mem[432] = 10'h16f;
        mem[433] = 10'h2b2;
        mem[434] = 10'h394;
        mem[435] = 10'h095;
        mem[436] = 10'h1b8;
        mem[437] = 10'h083;
        mem[438] = 10'h012;
        mem[439] = 10'h202;
        mem[440] = 10'h075;
        mem[441] = 10'h017;
        mem[442] = 10'h191;
        mem[443] = 10'h1bd;
        mem[444] = 10'h21f;
        mem[445] = 10'h1db;
        mem[446] = 10'h311;
        mem[447] = 10'h216;
        mem[448] = 10'h32e;
        mem[449] = 10'h1b7;
        mem[450] = 10'h057;
        mem[451] = 10'h361;
        mem[452] = 10'h331;
        mem[453] = 10'h362;
        mem[454] = 10'h2d4;
        mem[455] = 10'h1de;
        mem[456] = 10'h3e2;
        mem[457] = 10'h220;
        mem[458] = 10'h2f6;
        mem[459] = 10'h372;
        mem[460] = 10'h010;
        mem[461] = 10'h30a;
        mem[462] = 10'h051;
        mem[463] = 10'h310;
        mem[464] = 10'h320;
        mem[465] = 10'h325;
        mem[466] = 10'h0c3;
        mem[467] = 10'h3ef;
        mem[468] = 10'h2d9;
        mem[469] = 10'h1eb;
        mem[470] = 10'h143;
        mem[471] = 10'h0bb;
        mem[472] = 10'h0ca;
        mem[473] = 10'h3c5;
        mem[474] = 10'h24f;
        mem[475] = 10'h0dc;
        mem[476] = 10'h262;
        mem[477] = 10'h3cf;
        mem[478] = 10'h317;
        mem[479] = 10'h1c8;
        mem[480] = 10'h0fb;
        mem[481] = 10'h33c;
        mem[482] = 10'h172;
        mem[483] = 10'h3d8;
        mem[484] = 10'h388;
        mem[485] = 10'h25f;
        mem[486] = 10'h150;
        mem[487] = 10'h316;
        mem[488] = 10'h249;
        mem[489] = 10'h3d3;
        mem[490] = 10'h12a;
        mem[491] = 10'h1d5;
        mem[492] = 10'h233;
        mem[493] = 10'h274;
        mem[494] = 10'h27b;
        mem[495] = 10'h14c;
        mem[496] = 10'h09d;
        mem[497] = 10'h3de;
        mem[498] = 10'h387;
        mem[499] = 10'h33a;
        mem[500] = 10'h02a;
        mem[501] = 10'h013;
        mem[502] = 10'h1f4;
        mem[503] = 10'h276;
        mem[504] = 10'h23f;
        mem[505] = 10'h109;
        mem[506] = 10'h1b3;
        mem[507] = 10'h0fe;
        mem[508] = 10'h195;
        mem[509] = 10'h140;
        mem[510] = 10'h174;
        mem[511] = 10'h36a;
        mem[512] = 10'h24a;
        mem[513] = 10'h087;
        mem[514] = 10'h3d0;
        mem[515] = 10'h137;
        mem[516] = 10'h009;
        mem[517] = 10'h31b;
        mem[518] = 10'h227;
        mem[519] = 10'h17a;
        mem[520] = 10'h16c;
        mem[521] = 10'h17e;
        mem[522] = 10'h081;
        mem[523] = 10'h235;
        mem[524] = 10'h292;
        mem[525] = 10'h008;
        mem[526] = 10'h3bf;
        mem[527] = 10'h215;
        mem[528] = 10'h12e;
        mem[529] = 10'h24c;
        mem[530] = 10'h1b6;
        mem[531] = 10'h266;
        mem[532] = 10'h142;
        mem[533] = 10'h3ae;
        mem[534] = 10'h3ff;
        mem[535] = 10'h383;
        mem[536] = 10'h09e;
        mem[537] = 10'h01c;
        mem[538] = 10'h2b4;
        mem[539] = 10'h052;
        mem[540] = 10'h14b;
        mem[541] = 10'h3f2;
        mem[542] = 10'h33e;
        mem[543] = 10'h04b;
        mem[544] = 10'h342;
        mem[545] = 10'h1e9;
        mem[546] = 10'h3bb;
        mem[547] = 10'h13f;
        mem[548] = 10'h3c6;
        mem[549] = 10'h29e;
        mem[550] = 10'h182;
        mem[551] = 10'h028;
        mem[552] = 10'h1ff;
        mem[553] = 10'h1ed;
        mem[554] = 10'h3e7;
        mem[555] = 10'h315;
        mem[556] = 10'h299;
        mem[557] = 10'h34a;
        mem[558] = 10'h21b;
        mem[559] = 10'h3eb;
        mem[560] = 10'h099;
        mem[561] = 10'h14a;
        mem[562] = 10'h377;
        mem[563] = 10'h3b3;
        mem[564] = 10'h106;
        mem[565] = 10'h131;
        mem[566] = 10'h338;
        mem[567] = 10'h11b;
        mem[568] = 10'h3fe;
        mem[569] = 10'h2d8;
        mem[570] = 10'h357;
        mem[571] = 10'h072;
        mem[572] = 10'h3ce;
        mem[573] = 10'h0b4;
        mem[574] = 10'h32c;
        mem[575] = 10'h08a;
        mem[576] = 10'h2a3;
        mem[577] = 10'h037;
        mem[578] = 10'h035;
        mem[579] = 10'h21e;
        mem[580] = 10'h2a8;
        mem[581] = 10'h189;
        mem[582] = 10'h300;
        mem[583] = 10'h3fa;
        mem[584] = 10'h35e;
        mem[585] = 10'h34d;
        mem[586] = 10'h302;
        mem[587] = 10'h100;
        mem[588] = 10'h231;
        mem[589] = 10'h169;
        mem[590] = 10'h0ba;
        mem[591] = 10'h31e;
        mem[592] = 10'h0f6;
        mem[593] = 10'h00c;
        mem[594] = 10'h0e7;
        mem[595] = 10'h236;
        mem[596] = 10'h208;
        mem[597] = 10'h39a;
        mem[598] = 10'h1c3;
        mem[599] = 10'h159;
        mem[600] = 10'h1af;
        mem[601] = 10'h0db;
        mem[602] = 10'h1f9;
        mem[603] = 10'h05a;
        mem[604] = 10'h23d;
        mem[605] = 10'h264;
        mem[606] = 10'h35b;
        mem[607] = 10'h38f;
        mem[608] = 10'h282;
        mem[609] = 10'h024;
        mem[610] = 10'h38d;
        mem[611] = 10'h3a8;
        mem[612] = 10'h2cc;
        mem[613] = 10'h069;
        mem[614] = 10'h1b2;
        mem[615] = 10'h006;
        mem[616] = 10'h281;
        mem[617] = 10'h2fb;
        mem[618] = 10'h0f8;
        mem[619] = 10'h3ed;
        mem[620] = 10'h2d6;
        mem[621] = 10'h3bd;
        mem[622] = 10'h283;
        mem[623] = 10'h18b;
        mem[624] = 10'h2ee;
        mem[625] = 10'h322;
        mem[626] = 10'h2e6;
        mem[627] = 10'h323;
        mem[628] = 10'h391;
        mem[629] = 10'h181;
        mem[630] = 10'h288;
        mem[631] = 10'h04f;
        mem[632] = 10'h105;
        mem[633] = 10'h184;
        mem[634] = 10'h1f7;
        mem[635] = 10'h091;
        mem[636] = 10'h01b;
        mem[637] = 10'h1e5;
        mem[638] = 10'h118;
        mem[639] = 10'h170;
        mem[640] = 10'h0ec;
        mem[641] = 10'h01d;
        mem[642] = 10'h114;
        mem[643] = 10'h146;
        mem[644] = 10'h007;
        mem[645] = 10'h11c;
        mem[646] = 10'h152;
        mem[647] = 10'h2fa;
        mem[648] = 10'h02d;
        mem[649] = 10'h029;
        mem[650] = 10'h3f5;
        mem[651] = 10'h2da;
        mem[652] = 10'h3b5;
        mem[653] = 10'h2db;
        mem[654] = 10'h0e0;
        mem[655] = 10'h098;
        mem[656] = 10'h079;
        mem[657] = 10'h0f7;
        mem[658] = 10'h034;
        mem[659] = 10'h24b;
        mem[660] = 10'h12d;
        mem[661] = 10'h1fa;
        mem[662] = 10'h060;
        mem[663] = 10'h2aa;
        mem[664] = 10'h364;
        mem[665] = 10'h3db;
        mem[666] = 10'h036;
        mem[667] = 10'h1c2;
        mem[668] = 10'h019;
        mem[669] = 10'h244;
        mem[670] = 10'h15b;
        mem[671] = 10'h399;
        mem[672] = 10'h3ea;
        mem[673] = 10'h335;
        mem[674] = 10'h19c;
        mem[675] = 10'h0ed;
        mem[676] = 10'h2bb;
        mem[677] = 10'h148;
        mem[678] = 10'h3e4;
        mem[679] = 10'h3f6;
        mem[680] = 10'h379;
        mem[681] = 10'h0ab;
        mem[682] = 10'h273;
        mem[683] = 10'h126;
        mem[684] = 10'h267;
        mem[685] = 10'h294;
        mem[686] = 10'h0e5;
        mem[687] = 10'h003;
        mem[688] = 10'h270;
        mem[689] = 10'h15f;
        mem[690] = 10'h37c;
        mem[691] = 10'h329;
        mem[692] = 10'h03d;
        mem[693] = 10'h3f9;
        mem[694] = 10'h07a;
        mem[695] = 10'h192;
        mem[696] = 10'h055;
        mem[697] = 10'h018;
        mem[698] = 10'h068;
        mem[699] = 10'h1e4;
        mem[700] = 10'h1da;
        mem[701] = 10'h2f1;
        mem[702] = 10'h295;
        mem[703] = 10'h3b2;
        mem[704] = 10'h30d;
        mem[705] = 10'h290;
        mem[706] = 10'h3d6;
        mem[707] = 10'h111;
        mem[708] = 10'h0d7;
        mem[709] = 10'h026;
        mem[710] = 10'h2b1;
        mem[711] = 10'h065;
        mem[712] = 10'h02b;
        mem[713] = 10'h199;
        mem[714] = 10'h188;
        mem[715] = 10'h206;
        mem[716] = 10'h0ac;
        mem[717] = 10'h2e1;
        mem[718] = 10'h3cb;
        mem[719] = 10'h352;
        mem[720] = 10'h219;
        mem[721] = 10'h153;
        mem[722] = 10'h37d;
        mem[723] = 10'h06b;
        mem[724] = 10'h318;
        mem[725] = 10'h303;
        mem[726] = 10'h16e;
        mem[727] = 10'h09b;
        mem[728] = 10'h313;
        mem[729] = 10'h3e9;
        mem[730] = 10'h06e;
        mem[731] = 10'h375;
        mem[732] = 10'h393;
        mem[733] = 10'h10f;
        mem[734] = 10'h3c3;
        mem[735] = 10'h3d5;
        mem[736] = 10'h2e2;
        mem[737] = 10'h1e0;
        mem[738] = 10'h16a;
        mem[739] = 10'h3f3;
        mem[740] = 10'h256;
        mem[741] = 10'h36c;
        mem[742] = 10'h251;
        mem[743] = 10'h28b;
        mem[744] = 10'h08f;
        mem[745] = 10'h1c7;
        mem[746] = 10'h0d6;
        mem[747] = 10'h10e;
        mem[748] = 10'h1fb;
        mem[749] = 10'h337;
        mem[750] = 10'h0e9;
        mem[751] = 10'h194;
        mem[752] = 10'h046;
        mem[753] = 10'h25b;
        mem[754] = 10'h08c;
        mem[755] = 10'h23c;
        mem[756] = 10'h10a;
        mem[757] = 10'h3a1;
        mem[758] = 10'h2f9;
        mem[759] = 10'h1a7;
        mem[760] = 10'h25d;
        mem[761] = 10'h1ca;
        mem[762] = 10'h101;
        mem[763] = 10'h257;
        mem[764] = 10'h38b;
        mem[765] = 10'h3a6;
        mem[766] = 10'h0cd;
        mem[767] = 10'h247;
        mem[768] = 10'h06c;
        mem[769] = 10'h2bc;
        mem[770] = 10'h03e;
        mem[771] = 10'h3d4;
        mem[772] = 10'h04e;
        mem[773] = 10'h250;
        mem[774] = 10'h0be;
        mem[775] = 10'h355;
        mem[776] = 10'h01a;
        mem[777] = 10'h19b;
        mem[778] = 10'h245;
        mem[779] = 10'h1e1;
        mem[780] = 10'h2b8;
        mem[781] = 10'h26e;
        mem[782] = 10'h0b5;
        mem[783] = 10'h218;
        mem[784] = 10'h1d2;
        mem[785] = 10'h371;
        mem[786] = 10'h224;
        mem[787] = 10'h1bf;
        mem[788] = 10'h312;
        mem[789] = 10'h0a6;
        mem[790] = 10'h2c8;
        mem[791] = 10'h05f;
        mem[792] = 10'h197;
        mem[793] = 10'h0b9;
        mem[794] = 10'h243;
        mem[795] = 10'h226;
        mem[796] = 10'h23b;
        mem[797] = 10'h127;
        mem[798] = 10'h3a0;
        mem[799] = 10'h36f;
        mem[800] = 10'h32b;
        mem[801] = 10'h1fd;
        mem[802] = 10'h1cc;
        mem[803] = 10'h3df;
        mem[804] = 10'h158;
        mem[805] = 10'h067;
        mem[806] = 10'h3dd;
        mem[807] = 10'h2a1;
        mem[808] = 10'h175;
        mem[809] = 10'h3d7;
        mem[810] = 10'h26b;
        mem[811] = 10'h082;
        mem[812] = 10'h166;
        mem[813] = 10'h0cc;
        mem[814] = 10'h280;
        mem[815] = 10'h386;
        mem[816] = 10'h396;
        mem[817] = 10'h19d;
        mem[818] = 10'h0ef;
        mem[819] = 10'h070;
        mem[820] = 10'h0ad;
        mem[821] = 10'h3c7;
        mem[822] = 10'h07c;
        mem[823] = 10'h354;
        mem[824] = 10'h385;
        mem[825] = 10'h145;
        mem[826] = 10'h34e;
        mem[827] = 10'h0d9;
        mem[828] = 10'h0fd;
        mem[829] = 10'h3d2;
        mem[830] = 10'h144;
        mem[831] = 10'h356;
        mem[832] = 10'h08e;
        mem[833] = 10'h2ef;
        mem[834] = 10'h13d;
        mem[835] = 10'h16d;
        mem[836] = 10'h369;
        mem[837] = 10'h3ac;
        mem[838] = 10'h0cf;
        mem[839] = 10'h0df;
        mem[840] = 10'h1b5;
        mem[841] = 10'h25c;
        mem[842] = 10'h18e;
        mem[843] = 10'h1bb;
        mem[844] = 10'h2fc;
        mem[845] = 10'h254;
        mem[846] = 10'h011;
        mem[847] = 10'h2c0;
        mem[848] = 10'h2ad;
        mem[849] = 10'h0d5;
        mem[850] = 10'h2d2;
        mem[851] = 10'h1f3;
        mem[852] = 10'h2ca;
        mem[853] = 10'h22f;
        mem[854] = 10'h3fb;
        mem[855] = 10'h2be;
        mem[856] = 10'h0c0;
        mem[857] = 10'h35a;
        mem[858] = 10'h1ea;
        mem[859] = 10'h1cd;
        mem[860] = 10'h1cf;
        mem[861] = 10'h02e;
        mem[862] = 10'h24e;
        mem[863] = 10'h09c;
        mem[864] = 10'h33f;
        mem[865] = 10'h285;
        mem[866] = 10'h21c;
        mem[867] = 10'h38a;
        mem[868] = 10'h2c7;
        mem[869] = 10'h16b;
        mem[870] = 10'h05c;
        mem[871] = 10'h1e3;
        mem[872] = 10'h35c;
        mem[873] = 10'h327;
        mem[874] = 10'h171;
        mem[875] = 10'h063;
        mem[876] = 10'h21a;
        mem[877] = 10'h160;
        mem[878] = 10'h1c4;
        mem[879] = 10'h314;
        mem[880] = 10'h32f;
        mem[881] = 10'h133;
        mem[882] = 10'h033;
        mem[883] = 10'h308;
        mem[884] = 10'h15e;
        mem[885] = 10'h3b8;
        mem[886] = 10'h09a;
        mem[887] = 10'h390;
        mem[888] = 10'h10d;
        mem[889] = 10'h34c;
        mem[890] = 10'h225;
        mem[891] = 10'h289;
        mem[892] = 10'h344;
        mem[893] = 10'h28c;
        mem[894] = 10'h269;
        mem[895] = 10'h039;
        mem[896] = 10'h00d;
        mem[897] = 10'h324;
        mem[898] = 10'h389;
        mem[899] = 10'h027;
        mem[900] = 10'h0e8;
        mem[901] = 10'h2d5;
        mem[902] = 10'h1f0;
        mem[903] = 10'h113;
        mem[904] = 10'h0eb;
        mem[905] = 10'h3c0;
        mem[906] = 10'h2c5;
        mem[907] = 10'h1be;
        mem[908] = 10'h0e2;
        mem[909] = 10'h373;
        mem[910] = 10'h34b;
        mem[911] = 10'h07d;
        mem[912] = 10'h1aa;
        mem[913] = 10'h0f1;
        mem[914] = 10'h1a9;
        mem[915] = 10'h297;
        mem[916] = 10'h0aa;
        mem[917] = 10'h0bf;
        mem[918] = 10'h022;
        mem[919] = 10'h062;
        mem[920] = 10'h211;
        mem[921] = 10'h18a;
        mem[922] = 10'h054;
        mem[923] = 10'h1df;
        mem[924] = 10'h203;
        mem[925] = 10'h2c4;
        mem[926] = 10'h204;
        mem[927] = 10'h3b4;
        mem[928] = 10'h0c1;
        mem[929] = 10'h00b;
        mem[930] = 10'h12f;
        mem[931] = 10'h092;
        mem[932] = 10'h0c5;
        mem[933] = 10'h2d1;
        mem[934] = 10'h255;
        mem[935] = 10'h301;
        mem[936] = 10'h207;
        mem[937] = 10'h3a2;
        mem[938] = 10'h190;
        mem[939] = 10'h2a9;
        mem[940] = 10'h1c9;
        mem[941] = 10'h198;
        mem[942] = 10'h242;
        mem[943] = 10'h19e;
        mem[944] = 10'h284;
        mem[945] = 10'h1a3;
        mem[946] = 10'h047;
        mem[947] = 10'h11a;
        mem[948] = 10'h33b;
        mem[949] = 10'h13e;
        mem[950] = 10'h347;
        mem[951] = 10'h27a;
        mem[952] = 10'h246;
        mem[953] = 10'h2e4;
        mem[954] = 10'h29a;
        mem[955] = 10'h0b2;
        mem[956] = 10'h0a5;
        mem[957] = 10'h050;
        mem[958] = 10'h238;
        mem[959] = 10'h066;
        mem[960] = 10'h27c;
        mem[961] = 10'h367;
        mem[962] = 10'h333;
        mem[963] = 10'h0ea;
        mem[964] = 10'h279;
        mem[965] = 10'h17b;
        mem[966] = 10'h168;
        mem[967] = 10'h296;
        mem[968] = 10'h3af;
        mem[969] = 10'h004;
        mem[970] = 10'h3ca;
        mem[971] = 10'h15a;
        mem[972] = 10'h2af;
        mem[973] = 10'h1cb;
        mem[974] = 10'h180;
        mem[975] = 10'h36b;
        mem[976] = 10'h041;
        mem[977] = 10'h084;
        mem[978] = 10'h2b7;
        mem[979] = 10'h00e;
        mem[980] = 10'h077;
        mem[981] = 10'h26c;
        mem[982] = 10'h1a5;
        mem[983] = 10'h380;
        mem[984] = 10'h01e;
        mem[985] = 10'h3dc;
        mem[986] = 10'h336;
        mem[987] = 10'h186;
        mem[988] = 10'h1f2;
        mem[989] = 10'h1c1;
        mem[990] = 10'h2ce;
        mem[991] = 10'h1b1;
        mem[992] = 10'h27d;
        mem[993] = 10'h3bc;
        mem[994] = 10'h2a5;
        mem[995] = 10'h119;
        mem[996] = 10'h0b3;
        mem[997] = 10'h0f9;
        mem[998] = 10'h0e4;
        mem[999] = 10'h00f;
        mem[1000] = 10'h0fa;
        mem[1001] = 10'h0f3;
        mem[1002] = 10'h3e3;
        mem[1003] = 10'h2ea;
        mem[1004] = 10'h128;
        mem[1005] = 10'h125;
        mem[1006] = 10'h38e;
        mem[1007] = 10'h071;
        mem[1008] = 10'h252;
        mem[1009] = 10'h29b;
        mem[1010] = 10'h0a0;
        mem[1011] = 10'h3fc;
        mem[1012] = 10'h1a6;
        mem[1013] = 10'h185;
        mem[1014] = 10'h37f;
        mem[1015] = 10'h277;
        mem[1016] = 10'h110;
        mem[1017] = 10'h032;
        mem[1018] = 10'h108;
        mem[1019] = 10'h090;
        mem[1020] = 10'h2de;
        mem[1021] = 10'h048;
        mem[1022] = 10'h395;
        mem[1023] = 10'h129;
    end
endmodule

module encrypt_4apply_sboxes(clk, in, out);
    input clk;
    input [639:0] in;
    output [639:0] out;
    encrypt_4sbox_small0 sbox0inst(clk, in[5:0], out[5:0]);
    encrypt_4sbox_small1 sbox1inst(clk, in[21:16], out[21:16]);
    encrypt_4sbox_large0 sbox2inst(clk, in[15:6], in[31:22], out[15:6], out[31:22]);
    encrypt_4sbox_small2 sbox3inst(clk, in[37:32], out[37:32]);
    encrypt_4sbox_small3 sbox4inst(clk, in[53:48], out[53:48]);
    encrypt_4sbox_large0 sbox5inst(clk, in[47:38], in[63:54], out[47:38], out[63:54]);
    encrypt_4sbox_small4 sbox6inst(clk, in[69:64], out[69:64]);
    encrypt_4sbox_small5 sbox7inst(clk, in[85:80], out[85:80]);
    encrypt_4sbox_large1 sbox8inst(clk, in[79:70], in[95:86], out[79:70], out[95:86]);
    encrypt_4sbox_small6 sbox9inst(clk, in[101:96], out[101:96]);
    encrypt_4sbox_small7 sbox10inst(clk, in[117:112], out[117:112]);
    encrypt_4sbox_large1 sbox11inst(clk, in[111:102], in[127:118], out[111:102], out[127:118]);
    encrypt_4sbox_small8 sbox12inst(clk, in[133:128], out[133:128]);
    encrypt_4sbox_small9 sbox13inst(clk, in[149:144], out[149:144]);
    encrypt_4sbox_large2 sbox14inst(clk, in[143:134], in[159:150], out[143:134], out[159:150]);
    encrypt_4sbox_small10 sbox15inst(clk, in[165:160], out[165:160]);
    encrypt_4sbox_small11 sbox16inst(clk, in[181:176], out[181:176]);
    encrypt_4sbox_large2 sbox17inst(clk, in[175:166], in[191:182], out[175:166], out[191:182]);
    encrypt_4sbox_small12 sbox18inst(clk, in[197:192], out[197:192]);
    encrypt_4sbox_small13 sbox19inst(clk, in[213:208], out[213:208]);
    encrypt_4sbox_large3 sbox20inst(clk, in[207:198], in[223:214], out[207:198], out[223:214]);
    encrypt_4sbox_small14 sbox21inst(clk, in[229:224], out[229:224]);
    encrypt_4sbox_small15 sbox22inst(clk, in[245:240], out[245:240]);
    encrypt_4sbox_large3 sbox23inst(clk, in[239:230], in[255:246], out[239:230], out[255:246]);
    encrypt_4sbox_small16 sbox24inst(clk, in[261:256], out[261:256]);
    encrypt_4sbox_small17 sbox25inst(clk, in[277:272], out[277:272]);
    encrypt_4sbox_large4 sbox26inst(clk, in[271:262], in[287:278], out[271:262], out[287:278]);
    encrypt_4sbox_small18 sbox27inst(clk, in[293:288], out[293:288]);
    encrypt_4sbox_small19 sbox28inst(clk, in[309:304], out[309:304]);
    encrypt_4sbox_large4 sbox29inst(clk, in[303:294], in[319:310], out[303:294], out[319:310]);
    encrypt_4sbox_small20 sbox30inst(clk, in[325:320], out[325:320]);
    encrypt_4sbox_small21 sbox31inst(clk, in[341:336], out[341:336]);
    encrypt_4sbox_large5 sbox32inst(clk, in[335:326], in[351:342], out[335:326], out[351:342]);
    encrypt_4sbox_small22 sbox33inst(clk, in[357:352], out[357:352]);
    encrypt_4sbox_small23 sbox34inst(clk, in[373:368], out[373:368]);
    encrypt_4sbox_large5 sbox35inst(clk, in[367:358], in[383:374], out[367:358], out[383:374]);
    encrypt_4sbox_small24 sbox36inst(clk, in[389:384], out[389:384]);
    encrypt_4sbox_small25 sbox37inst(clk, in[405:400], out[405:400]);
    encrypt_4sbox_large6 sbox38inst(clk, in[399:390], in[415:406], out[399:390], out[415:406]);
    encrypt_4sbox_small26 sbox39inst(clk, in[421:416], out[421:416]);
    encrypt_4sbox_small27 sbox40inst(clk, in[437:432], out[437:432]);
    encrypt_4sbox_large6 sbox41inst(clk, in[431:422], in[447:438], out[431:422], out[447:438]);
    encrypt_4sbox_small28 sbox42inst(clk, in[453:448], out[453:448]);
    encrypt_4sbox_small29 sbox43inst(clk, in[469:464], out[469:464]);
    encrypt_4sbox_large7 sbox44inst(clk, in[463:454], in[479:470], out[463:454], out[479:470]);
    encrypt_4sbox_small30 sbox45inst(clk, in[485:480], out[485:480]);
    encrypt_4sbox_small31 sbox46inst(clk, in[501:496], out[501:496]);
    encrypt_4sbox_large7 sbox47inst(clk, in[495:486], in[511:502], out[495:486], out[511:502]);
    encrypt_4sbox_small32 sbox48inst(clk, in[517:512], out[517:512]);
    encrypt_4sbox_small33 sbox49inst(clk, in[533:528], out[533:528]);
    encrypt_4sbox_large8 sbox50inst(clk, in[527:518], in[543:534], out[527:518], out[543:534]);
    encrypt_4sbox_small34 sbox51inst(clk, in[549:544], out[549:544]);
    encrypt_4sbox_small35 sbox52inst(clk, in[565:560], out[565:560]);
    encrypt_4sbox_large8 sbox53inst(clk, in[559:550], in[575:566], out[559:550], out[575:566]);
    encrypt_4sbox_small36 sbox54inst(clk, in[581:576], out[581:576]);
    encrypt_4sbox_small37 sbox55inst(clk, in[597:592], out[597:592]);
    encrypt_4sbox_large9 sbox56inst(clk, in[591:582], in[607:598], out[591:582], out[607:598]);
    encrypt_4sbox_small38 sbox57inst(clk, in[613:608], out[613:608]);
    encrypt_4sbox_small39 sbox58inst(clk, in[629:624], out[629:624]);
    encrypt_4sbox_large9 sbox59inst(clk, in[623:614], in[639:630], out[623:614], out[639:630]);
endmodule

module encrypt_4apply_pbox0(in, out);
    input [639:0] in;
    output [639:0] out;
    assign out[339] = in[0];
    assign out[287] = in[1];
    assign out[22] = in[2];
    assign out[521] = in[3];
    assign out[279] = in[4];
    assign out[371] = in[5];
    assign out[37] = in[6];
    assign out[540] = in[7];
    assign out[504] = in[8];
    assign out[308] = in[9];
    assign out[506] = in[10];
    assign out[310] = in[11];
    assign out[151] = in[12];
    assign out[525] = in[13];
    assign out[385] = in[14];
    assign out[110] = in[15];
    assign out[184] = in[16];
    assign out[388] = in[17];
    assign out[453] = in[18];
    assign out[119] = in[19];
    assign out[13] = in[20];
    assign out[307] = in[21];
    assign out[411] = in[22];
    assign out[288] = in[23];
    assign out[553] = in[24];
    assign out[618] = in[25];
    assign out[557] = in[26];
    assign out[482] = in[27];
    assign out[463] = in[28];
    assign out[501] = in[29];
    assign out[359] = in[30];
    assign out[269] = in[31];
    assign out[127] = in[32];
    assign out[488] = in[33];
    assign out[67] = in[34];
    assign out[163] = in[35];
    assign out[365] = in[36];
    assign out[366] = in[37];
    assign out[631] = in[38];
    assign out[378] = in[39];
    assign out[571] = in[40];
    assign out[102] = in[41];
    assign out[410] = in[42];
    assign out[150] = in[43];
    assign out[577] = in[44];
    assign out[12] = in[45];
    assign out[200] = in[46];
    assign out[239] = in[47];
    assign out[81] = in[48];
    assign out[440] = in[49];
    assign out[272] = in[50];
    assign out[419] = in[51];
    assign out[223] = in[52];
    assign out[328] = in[53];
    assign out[111] = in[54];
    assign out[48] = in[55];
    assign out[6] = in[56];
    assign out[93] = in[57];
    assign out[94] = in[58];
    assign out[513] = in[59];
    assign out[346] = in[60];
    assign out[283] = in[61];
    assign out[591] = in[62];
    assign out[60] = in[63];
    assign out[389] = in[64];
    assign out[330] = in[65];
    assign out[123] = in[66];
    assign out[456] = in[67];
    assign out[348] = in[68];
    assign out[144] = in[69];
    assign out[539] = in[70];
    assign out[437] = in[71];
    assign out[507] = in[72];
    assign out[517] = in[73];
    assign out[46] = in[74];
    assign out[108] = in[75];
    assign out[530] = in[76];
    assign out[421] = in[77];
    assign out[71] = in[78];
    assign out[143] = in[79];
    assign out[212] = in[80];
    assign out[220] = in[81];
    assign out[551] = in[82];
    assign out[158] = in[83];
    assign out[592] = in[84];
    assign out[18] = in[85];
    assign out[361] = in[86];
    assign out[531] = in[87];
    assign out[392] = in[88];
    assign out[221] = in[89];
    assign out[301] = in[90];
    assign out[599] = in[91];
    assign out[623] = in[92];
    assign out[420] = in[93];
    assign out[63] = in[94];
    assign out[92] = in[95];
    assign out[629] = in[96];
    assign out[626] = in[97];
    assign out[112] = in[98];
    assign out[257] = in[99];
    assign out[72] = in[100];
    assign out[197] = in[101];
    assign out[99] = in[102];
    assign out[615] = in[103];
    assign out[475] = in[104];
    assign out[201] = in[105];
    assign out[472] = in[106];
    assign out[576] = in[107];
    assign out[11] = in[108];
    assign out[59] = in[109];
    assign out[79] = in[110];
    assign out[512] = in[111];
    assign out[624] = in[112];
    assign out[69] = in[113];
    assign out[441] = in[114];
    assign out[395] = in[115];
    assign out[583] = in[116];
    assign out[382] = in[117];
    assign out[74] = in[118];
    assign out[563] = in[119];
    assign out[422] = in[120];
    assign out[384] = in[121];
    assign out[323] = in[122];
    assign out[187] = in[123];
    assign out[121] = in[124];
    assign out[360] = in[125];
    assign out[216] = in[126];
    assign out[493] = in[127];
    assign out[254] = in[128];
    assign out[397] = in[129];
    assign out[496] = in[130];
    assign out[253] = in[131];
    assign out[50] = in[132];
    assign out[115] = in[133];
    assign out[625] = in[134];
    assign out[122] = in[135];
    assign out[502] = in[136];
    assign out[390] = in[137];
    assign out[565] = in[138];
    assign out[148] = in[139];
    assign out[275] = in[140];
    assign out[0] = in[141];
    assign out[267] = in[142];
    assign out[569] = in[143];
    assign out[149] = in[144];
    assign out[276] = in[145];
    assign out[9] = in[146];
    assign out[316] = in[147];
    assign out[217] = in[148];
    assign out[218] = in[149];
    assign out[473] = in[150];
    assign out[350] = in[151];
    assign out[321] = in[152];
    assign out[548] = in[153];
    assign out[344] = in[154];
    assign out[73] = in[155];
    assign out[519] = in[156];
    assign out[157] = in[157];
    assign out[227] = in[158];
    assign out[560] = in[159];
    assign out[555] = in[160];
    assign out[523] = in[161];
    assign out[10] = in[162];
    assign out[564] = in[163];
    assign out[487] = in[164];
    assign out[170] = in[165];
    assign out[20] = in[166];
    assign out[405] = in[167];
    assign out[232] = in[168];
    assign out[87] = in[169];
    assign out[168] = in[170];
    assign out[429] = in[171];
    assign out[298] = in[172];
    assign out[38] = in[173];
    assign out[238] = in[174];
    assign out[425] = in[175];
    assign out[30] = in[176];
    assign out[633] = in[177];
    assign out[373] = in[178];
    assign out[542] = in[179];
    assign out[39] = in[180];
    assign out[518] = in[181];
    assign out[484] = in[182];
    assign out[514] = in[183];
    assign out[536] = in[184];
    assign out[586] = in[185];
    assign out[538] = in[186];
    assign out[41] = in[187];
    assign out[614] = in[188];
    assign out[457] = in[189];
    assign out[53] = in[190];
    assign out[381] = in[191];
    assign out[619] = in[192];
    assign out[510] = in[193];
    assign out[106] = in[194];
    assign out[621] = in[195];
    assign out[559] = in[196];
    assign out[447] = in[197];
    assign out[393] = in[198];
    assign out[270] = in[199];
    assign out[247] = in[200];
    assign out[327] = in[201];
    assign out[461] = in[202];
    assign out[3] = in[203];
    assign out[116] = in[204];
    assign out[141] = in[205];
    assign out[7] = in[206];
    assign out[137] = in[207];
    assign out[202] = in[208];
    assign out[203] = in[209];
    assign out[277] = in[210];
    assign out[130] = in[211];
    assign out[142] = in[212];
    assign out[407] = in[213];
    assign out[349] = in[214];
    assign out[198] = in[215];
    assign out[17] = in[216];
    assign out[459] = in[217];
    assign out[476] = in[218];
    assign out[224] = in[219];
    assign out[83] = in[220];
    assign out[16] = in[221];
    assign out[21] = in[222];
    assign out[228] = in[223];
    assign out[492] = in[224];
    assign out[155] = in[225];
    assign out[297] = in[226];
    assign out[469] = in[227];
    assign out[354] = in[228];
    assign out[630] = in[229];
    assign out[434] = in[230];
    assign out[236] = in[231];
    assign out[584] = in[232];
    assign out[152] = in[233];
    assign out[562] = in[234];
    assign out[176] = in[235];
    assign out[494] = in[236];
    assign out[27] = in[237];
    assign out[491] = in[238];
    assign out[169] = in[239];
    assign out[508] = in[240];
    assign out[436] = in[241];
    assign out[579] = in[242];
    assign out[314] = in[243];
    assign out[109] = in[244];
    assign out[312] = in[245];
    assign out[450] = in[246];
    assign out[47] = in[247];
    assign out[248] = in[248];
    assign out[612] = in[249];
    assign out[250] = in[250];
    assign out[128] = in[251];
    assign out[182] = in[252];
    assign out[511] = in[253];
    assign out[55] = in[254];
    assign out[262] = in[255];
    assign out[320] = in[256];
    assign out[529] = in[257];
    assign out[258] = in[258];
    assign out[467] = in[259];
    assign out[164] = in[260];
    assign out[80] = in[261];
    assign out[580] = in[262];
    assign out[125] = in[263];
    assign out[460] = in[264];
    assign out[209] = in[265];
    assign out[135] = in[266];
    assign out[140] = in[267];
    assign out[205] = in[268];
    assign out[89] = in[269];
    assign out[544] = in[270];
    assign out[477] = in[271];
    assign out[402] = in[272];
    assign out[337] = in[273];
    assign out[107] = in[274];
    assign out[547] = in[275];
    assign out[180] = in[276];
    assign out[146] = in[277];
    assign out[278] = in[278];
    assign out[34] = in[279];
    assign out[100] = in[280];
    assign out[19] = in[281];
    assign out[535] = in[282];
    assign out[292] = in[283];
    assign out[244] = in[284];
    assign out[40] = in[285];
    assign out[84] = in[286];
    assign out[43] = in[287];
    assign out[86] = in[288];
    assign out[226] = in[289];
    assign out[266] = in[290];
    assign out[464] = in[291];
    assign out[225] = in[292];
    assign out[91] = in[293];
    assign out[500] = in[294];
    assign out[33] = in[295];
    assign out[596] = in[296];
    assign out[35] = in[297];
    assign out[274] = in[298];
    assign out[194] = in[299];
    assign out[430] = in[300];
    assign out[120] = in[301];
    assign out[432] = in[302];
    assign out[497] = in[303];
    assign out[173] = in[304];
    assign out[145] = in[305];
    assign out[179] = in[306];
    assign out[329] = in[307];
    assign out[246] = in[308];
    assign out[439] = in[309];
    assign out[546] = in[310];
    assign out[113] = in[311];
    assign out[454] = in[312];
    assign out[153] = in[313];
    assign out[516] = in[314];
    assign out[189] = in[315];
    assign out[570] = in[316];
    assign out[326] = in[317];
    assign out[222] = in[318];
    assign out[88] = in[319];
    assign out[594] = in[320];
    assign out[131] = in[321];
    assign out[264] = in[322];
    assign out[132] = in[323];
    assign out[62] = in[324];
    assign out[229] = in[325];
    assign out[458] = in[326];
    assign out[336] = in[327];
    assign out[452] = in[328];
    assign out[139] = in[329];
    assign out[408] = in[330];
    assign out[342] = in[331];
    assign out[522] = in[332];
    assign out[401] = in[333];
    assign out[600] = in[334];
    assign out[609] = in[335];
    assign out[210] = in[336];
    assign out[28] = in[337];
    assign out[211] = in[338];
    assign out[605] = in[339];
    assign out[593] = in[340];
    assign out[607] = in[341];
    assign out[299] = in[342];
    assign out[403] = in[343];
    assign out[213] = in[344];
    assign out[154] = in[345];
    assign out[304] = in[346];
    assign out[415] = in[347];
    assign out[478] = in[348];
    assign out[54] = in[349];
    assign out[474] = in[350];
    assign out[42] = in[351];
    assign out[192] = in[352];
    assign out[249] = in[353];
    assign out[590] = in[354];
    assign out[195] = in[355];
    assign out[480] = in[356];
    assign out[31] = in[357];
    assign out[231] = in[358];
    assign out[549] = in[359];
    assign out[255] = in[360];
    assign out[230] = in[361];
    assign out[534] = in[362];
    assign out[68] = in[363];
    assign out[196] = in[364];
    assign out[70] = in[365];
    assign out[313] = in[366];
    assign out[325] = in[367];
    assign out[604] = in[368];
    assign out[435] = in[369];
    assign out[370] = in[370];
    assign out[240] = in[371];
    assign out[481] = in[372];
    assign out[65] = in[373];
    assign out[331] = in[374];
    assign out[322] = in[375];
    assign out[185] = in[376];
    assign out[509] = in[377];
    assign out[271] = in[378];
    assign out[355] = in[379];
    assign out[114] = in[380];
    assign out[527] = in[381];
    assign out[191] = in[382];
    assign out[199] = in[383];
    assign out[204] = in[384];
    assign out[256] = in[385];
    assign out[455] = in[386];
    assign out[36] = in[387];
    assign out[101] = in[388];
    assign out[380] = in[389];
    assign out[515] = in[390];
    assign out[442] = in[391];
    assign out[396] = in[392];
    assign out[25] = in[393];
    assign out[85] = in[394];
    assign out[637] = in[395];
    assign out[574] = in[396];
    assign out[268] = in[397];
    assign out[64] = in[398];
    assign out[95] = in[399];
    assign out[332] = in[400];
    assign out[628] = in[401];
    assign out[406] = in[402];
    assign out[532] = in[403];
    assign out[188] = in[404];
    assign out[568] = in[405];
    assign out[338] = in[406];
    assign out[8] = in[407];
    assign out[601] = in[408];
    assign out[280] = in[409];
    assign out[166] = in[410];
    assign out[347] = in[411];
    assign out[294] = in[412];
    assign out[177] = in[413];
    assign out[528] = in[414];
    assign out[351] = in[415];
    assign out[352] = in[416];
    assign out[44] = in[417];
    assign out[219] = in[418];
    assign out[423] = in[419];
    assign out[387] = in[420];
    assign out[241] = in[421];
    assign out[159] = in[422];
    assign out[427] = in[423];
    assign out[295] = in[424];
    assign out[259] = in[425];
    assign out[117] = in[426];
    assign out[362] = in[427];
    assign out[291] = in[428];
    assign out[78] = in[429];
    assign out[57] = in[430];
    assign out[377] = in[431];
    assign out[483] = in[432];
    assign out[175] = in[433];
    assign out[61] = in[434];
    assign out[556] = in[435];
    assign out[1] = in[436];
    assign out[305] = in[437];
    assign out[400] = in[438];
    assign out[273] = in[439];
    assign out[311] = in[440];
    assign out[208] = in[441];
    assign out[134] = in[442];
    assign out[448] = in[443];
    assign out[245] = in[444];
    assign out[613] = in[445];
    assign out[567] = in[446];
    assign out[318] = in[447];
    assign out[375] = in[448];
    assign out[428] = in[449];
    assign out[412] = in[450];
    assign out[333] = in[451];
    assign out[15] = in[452];
    assign out[156] = in[453];
    assign out[575] = in[454];
    assign out[289] = in[455];
    assign out[58] = in[456];
    assign out[398] = in[457];
    assign out[242] = in[458];
    assign out[124] = in[459];
    assign out[45] = in[460];
    assign out[526] = in[461];
    assign out[14] = in[462];
    assign out[386] = in[463];
    assign out[426] = in[464];
    assign out[363] = in[465];
    assign out[566] = in[466];
    assign out[96] = in[467];
    assign out[302] = in[468];
    assign out[573] = in[469];
    assign out[638] = in[470];
    assign out[369] = in[471];
    assign out[104] = in[472];
    assign out[414] = in[473];
    assign out[479] = in[474];
    assign out[282] = in[475];
    assign out[639] = in[476];
    assign out[281] = in[477];
    assign out[286] = in[478];
    assign out[446] = in[479];
    assign out[520] = in[480];
    assign out[285] = in[481];
    assign out[486] = in[482];
    assign out[424] = in[483];
    assign out[162] = in[484];
    assign out[550] = in[485];
    assign out[186] = in[486];
    assign out[165] = in[487];
    assign out[524] = in[488];
    assign out[90] = in[489];
    assign out[353] = in[490];
    assign out[29] = in[491];
    assign out[374] = in[492];
    assign out[300] = in[493];
    assign out[167] = in[494];
    assign out[552] = in[495];
    assign out[367] = in[496];
    assign out[136] = in[497];
    assign out[485] = in[498];
    assign out[503] = in[499];
    assign out[237] = in[500];
    assign out[319] = in[501];
    assign out[23] = in[502];
    assign out[603] = in[503];
    assign out[561] = in[504];
    assign out[634] = in[505];
    assign out[541] = in[506];
    assign out[75] = in[507];
    assign out[622] = in[508];
    assign out[545] = in[509];
    assign out[317] = in[510];
    assign out[379] = in[511];
    assign out[433] = in[512];
    assign out[252] = in[513];
    assign out[611] = in[514];
    assign out[190] = in[515];
    assign out[589] = in[516];
    assign out[52] = in[517];
    assign out[2] = in[518];
    assign out[118] = in[519];
    assign out[505] = in[520];
    assign out[133] = in[521];
    assign out[616] = in[522];
    assign out[602] = in[523];
    assign out[376] = in[524];
    assign out[315] = in[525];
    assign out[620] = in[526];
    assign out[138] = in[527];
    assign out[5] = in[528];
    assign out[383] = in[529];
    assign out[343] = in[530];
    assign out[610] = in[531];
    assign out[399] = in[532];
    assign out[627] = in[533];
    assign out[471] = in[534];
    assign out[76] = in[535];
    assign out[4] = in[536];
    assign out[404] = in[537];
    assign out[635] = in[538];
    assign out[263] = in[539];
    assign out[413] = in[540];
    assign out[260] = in[541];
    assign out[636] = in[542];
    assign out[466] = in[543];
    assign out[465] = in[544];
    assign out[126] = in[545];
    assign out[449] = in[546];
    assign out[468] = in[547];
    assign out[578] = in[548];
    assign out[558] = in[549];
    assign out[98] = in[550];
    assign out[234] = in[551];
    assign out[335] = in[552];
    assign out[26] = in[553];
    assign out[303] = in[554];
    assign out[174] = in[555];
    assign out[24] = in[556];
    assign out[409] = in[557];
    assign out[495] = in[558];
    assign out[235] = in[559];
    assign out[171] = in[560];
    assign out[214] = in[561];
    assign out[595] = in[562];
    assign out[364] = in[563];
    assign out[32] = in[564];
    assign out[82] = in[565];
    assign out[418] = in[566];
    assign out[470] = in[567];
    assign out[105] = in[568];
    assign out[357] = in[569];
    assign out[193] = in[570];
    assign out[372] = in[571];
    assign out[161] = in[572];
    assign out[554] = in[573];
    assign out[490] = in[574];
    assign out[608] = in[575];
    assign out[585] = in[576];
    assign out[444] = in[577];
    assign out[51] = in[578];
    assign out[56] = in[579];
    assign out[97] = in[580];
    assign out[129] = in[581];
    assign out[391] = in[582];
    assign out[499] = in[583];
    assign out[451] = in[584];
    assign out[309] = in[585];
    assign out[103] = in[586];
    assign out[632] = in[587];
    assign out[533] = in[588];
    assign out[598] = in[589];
    assign out[243] = in[590];
    assign out[606] = in[591];
    assign out[543] = in[592];
    assign out[445] = in[593];
    assign out[183] = in[594];
    assign out[66] = in[595];
    assign out[49] = in[596];
    assign out[334] = in[597];
    assign out[251] = in[598];
    assign out[261] = in[599];
    assign out[147] = in[600];
    assign out[394] = in[601];
    assign out[341] = in[602];
    assign out[215] = in[603];
    assign out[443] = in[604];
    assign out[160] = in[605];
    assign out[77] = in[606];
    assign out[356] = in[607];
    assign out[617] = in[608];
    assign out[284] = in[609];
    assign out[265] = in[610];
    assign out[296] = in[611];
    assign out[581] = in[612];
    assign out[582] = in[613];
    assign out[417] = in[614];
    assign out[290] = in[615];
    assign out[340] = in[616];
    assign out[206] = in[617];
    assign out[207] = in[618];
    assign out[178] = in[619];
    assign out[293] = in[620];
    assign out[416] = in[621];
    assign out[233] = in[622];
    assign out[462] = in[623];
    assign out[172] = in[624];
    assign out[498] = in[625];
    assign out[345] = in[626];
    assign out[572] = in[627];
    assign out[597] = in[628];
    assign out[368] = in[629];
    assign out[489] = in[630];
    assign out[306] = in[631];
    assign out[537] = in[632];
    assign out[181] = in[633];
    assign out[358] = in[634];
    assign out[438] = in[635];
    assign out[587] = in[636];
    assign out[588] = in[637];
    assign out[431] = in[638];
    assign out[324] = in[639];
endmodule

module encrypt_4apply_pbox1(in, out);
    input [639:0] in;
    output [639:0] out;
    assign out[244] = in[0];
    assign out[414] = in[1];
    assign out[466] = in[2];
    assign out[50] = in[3];
    assign out[220] = in[4];
    assign out[405] = in[5];
    assign out[186] = in[6];
    assign out[575] = in[7];
    assign out[397] = in[8];
    assign out[574] = in[9];
    assign out[113] = in[10];
    assign out[424] = in[11];
    assign out[588] = in[12];
    assign out[589] = in[13];
    assign out[346] = in[14];
    assign out[516] = in[15];
    assign out[232] = in[16];
    assign out[290] = in[17];
    assign out[434] = in[18];
    assign out[419] = in[19];
    assign out[524] = in[20];
    assign out[485] = in[21];
    assign out[62] = in[22];
    assign out[291] = in[23];
    assign out[271] = in[24];
    assign out[300] = in[25];
    assign out[273] = in[26];
    assign out[218] = in[27];
    assign out[532] = in[28];
    assign out[209] = in[29];
    assign out[369] = in[30];
    assign out[583] = in[31];
    assign out[184] = in[32];
    assign out[282] = in[33];
    assign out[74] = in[34];
    assign out[163] = in[35];
    assign out[449] = in[36];
    assign out[240] = in[37];
    assign out[85] = in[38];
    assign out[607] = in[39];
    assign out[545] = in[40];
    assign out[609] = in[41];
    assign out[374] = in[42];
    assign out[555] = in[43];
    assign out[613] = in[44];
    assign out[493] = in[45];
    assign out[550] = in[46];
    assign out[87] = in[47];
    assign out[600] = in[48];
    assign out[252] = in[49];
    assign out[299] = in[50];
    assign out[383] = in[51];
    assign out[243] = in[52];
    assign out[29] = in[53];
    assign out[454] = in[54];
    assign out[31] = in[55];
    assign out[32] = in[56];
    assign out[304] = in[57];
    assign out[506] = in[58];
    assign out[395] = in[59];
    assign out[344] = in[60];
    assign out[310] = in[61];
    assign out[375] = in[62];
    assign out[217] = in[63];
    assign out[631] = in[64];
    assign out[553] = in[65];
    assign out[142] = in[66];
    assign out[43] = in[67];
    assign out[343] = in[68];
    assign out[45] = in[69];
    assign out[338] = in[70];
    assign out[519] = in[71];
    assign out[135] = in[72];
    assign out[512] = in[73];
    assign out[347] = in[74];
    assign out[411] = in[75];
    assign out[140] = in[76];
    assign out[167] = in[77];
    assign out[491] = in[78];
    assign out[479] = in[79];
    assign out[120] = in[80];
    assign out[56] = in[81];
    assign out[109] = in[82];
    assign out[123] = in[83];
    assign out[420] = in[84];
    assign out[526] = in[85];
    assign out[161] = in[86];
    assign out[296] = in[87];
    assign out[593] = in[88];
    assign out[116] = in[89];
    assign out[66] = in[90];
    assign out[181] = in[91];
    assign out[155] = in[92];
    assign out[377] = in[93];
    assign out[518] = in[94];
    assign out[7] = in[95];
    assign out[212] = in[96];
    assign out[317] = in[97];
    assign out[72] = in[98];
    assign out[547] = in[99];
    assign out[283] = in[100];
    assign out[541] = in[101];
    assign out[543] = in[102];
    assign out[439] = in[103];
    assign out[287] = in[104];
    assign out[4] = in[105];
    assign out[455] = in[106];
    assign out[456] = in[107];
    assign out[620] = in[108];
    assign out[185] = in[109];
    assign out[598] = in[110];
    assign out[358] = in[111];
    assign out[164] = in[112];
    assign out[462] = in[113];
    assign out[318] = in[114];
    assign out[27] = in[115];
    assign out[327] = in[116];
    assign out[437] = in[117];
    assign out[144] = in[118];
    assign out[339] = in[119];
    assign out[392] = in[120];
    assign out[330] = in[121];
    assign out[474] = in[122];
    assign out[627] = in[123];
    assign out[36] = in[124];
    assign out[24] = in[125];
    assign out[25] = in[126];
    assign out[615] = in[127];
    assign out[503] = in[128];
    assign out[406] = in[129];
    assign out[214] = in[130];
    assign out[54] = in[131];
    assign out[604] = in[132];
    assign out[410] = in[133];
    assign out[157] = in[134];
    assign out[219] = in[135];
    assign out[584] = in[136];
    assign out[448] = in[137];
    assign out[222] = in[138];
    assign out[334] = in[139];
    assign out[224] = in[140];
    assign out[191] = in[141];
    assign out[435] = in[142];
    assign out[569] = in[143];
    assign out[0] = in[144];
    assign out[635] = in[145];
    assign out[393] = in[146];
    assign out[280] = in[147];
    assign out[556] = in[148];
    assign out[89] = in[149];
    assign out[576] = in[150];
    assign out[471] = in[151];
    assign out[408] = in[152];
    assign out[12] = in[153];
    assign out[128] = in[154];
    assign out[380] = in[155];
    assign out[497] = in[156];
    assign out[207] = in[157];
    assign out[17] = in[158];
    assign out[197] = in[159];
    assign out[146] = in[160];
    assign out[276] = in[161];
    assign out[614] = in[162];
    assign out[342] = in[163];
    assign out[636] = in[164];
    assign out[637] = in[165];
    assign out[263] = in[166];
    assign out[572] = in[167];
    assign out[509] = in[168];
    assign out[192] = in[169];
    assign out[46] = in[170];
    assign out[332] = in[171];
    assign out[385] = in[172];
    assign out[450] = in[173];
    assign out[335] = in[174];
    assign out[580] = in[175];
    assign out[150] = in[176];
    assign out[622] = in[177];
    assign out[391] = in[178];
    assign out[475] = in[179];
    assign out[628] = in[180];
    assign out[101] = in[181];
    assign out[587] = in[182];
    assign out[494] = in[183];
    assign out[528] = in[184];
    assign out[108] = in[185];
    assign out[527] = in[186];
    assign out[160] = in[187];
    assign out[481] = in[188];
    assign out[594] = in[189];
    assign out[467] = in[190];
    assign out[579] = in[191];
    assign out[353] = in[192];
    assign out[52] = in[193];
    assign out[70] = in[194];
    assign out[536] = in[195];
    assign out[601] = in[196];
    assign out[376] = in[197];
    assign out[329] = in[198];
    assign out[409] = in[199];
    assign out[156] = in[200];
    assign out[124] = in[201];
    assign out[415] = in[202];
    assign out[608] = in[203];
    assign out[63] = in[204];
    assign out[256] = in[205];
    assign out[483] = in[206];
    assign out[2] = in[207];
    assign out[84] = in[208];
    assign out[370] = in[209];
    assign out[371] = in[210];
    assign out[308] = in[211];
    assign out[459] = in[212];
    assign out[233] = in[213];
    assign out[173] = in[214];
    assign out[425] = in[215];
    assign out[426] = in[216];
    assign out[558] = in[217];
    assign out[623] = in[218];
    assign out[560] = in[219];
    assign out[625] = in[220];
    assign out[389] = in[221];
    assign out[178] = in[222];
    assign out[18] = in[223];
    assign out[480] = in[224];
    assign out[523] = in[225];
    assign out[48] = in[226];
    assign out[360] = in[227];
    assign out[361] = in[228];
    assign out[591] = in[229];
    assign out[204] = in[230];
    assign out[26] = in[231];
    assign out[188] = in[232];
    assign out[446] = in[233];
    assign out[93] = in[234];
    assign out[403] = in[235];
    assign out[492] = in[236];
    assign out[96] = in[237];
    assign out[30] = in[238];
    assign out[559] = in[239];
    assign out[564] = in[240];
    assign out[585] = in[241];
    assign out[134] = in[242];
    assign out[229] = in[243];
    assign out[561] = in[244];
    assign out[154] = in[245];
    assign out[41] = in[246];
    assign out[42] = in[247];
    assign out[394] = in[248];
    assign out[432] = in[249];
    assign out[418] = in[250];
    assign out[549] = in[251];
    assign out[401] = in[252];
    assign out[321] = in[253];
    assign out[322] = in[254];
    assign out[596] = in[255];
    assign out[307] = in[256];
    assign out[624] = in[257];
    assign out[176] = in[258];
    assign out[226] = in[259];
    assign out[387] = in[260];
    assign out[179] = in[261];
    assign out[490] = in[262];
    assign out[129] = in[263];
    assign out[246] = in[264];
    assign out[131] = in[265];
    assign out[573] = in[266];
    assign out[5] = in[267];
    assign out[71] = in[268];
    assign out[249] = in[269];
    assign out[9] = in[270];
    assign out[238] = in[271];
    assign out[487] = in[272];
    assign out[464] = in[273];
    assign out[567] = in[274];
    assign out[429] = in[275];
    assign out[79] = in[276];
    assign out[505] = in[277];
    assign out[132] = in[278];
    assign out[266] = in[279];
    assign out[570] = in[280];
    assign out[211] = in[281];
    assign out[187] = in[282];
    assign out[44] = in[283];
    assign out[114] = in[284];
    assign out[254] = in[285];
    assign out[253] = in[286];
    assign out[513] = in[287];
    assign out[193] = in[288];
    assign out[453] = in[289];
    assign out[597] = in[290];
    assign out[143] = in[291];
    assign out[443] = in[292];
    assign out[223] = in[293];
    assign out[345] = in[294];
    assign out[537] = in[295];
    assign out[423] = in[296];
    assign out[348] = in[297];
    assign out[489] = in[298];
    assign out[255] = in[299];
    assign out[441] = in[300];
    assign out[388] = in[301];
    assign out[284] = in[302];
    assign out[546] = in[303];
    assign out[404] = in[304];
    assign out[316] = in[305];
    assign out[172] = in[306];
    assign out[498] = in[307];
    assign out[639] = in[308];
    assign out[227] = in[309];
    assign out[356] = in[310];
    assign out[465] = in[311];
    assign out[73] = in[312];
    assign out[313] = in[313];
    assign out[557] = in[314];
    assign out[363] = in[315];
    assign out[77] = in[316];
    assign out[328] = in[317];
    assign out[170] = in[318];
    assign out[522] = in[319];
    assign out[81] = in[320];
    assign out[162] = in[321];
    assign out[333] = in[322];
    assign out[336] = in[323];
    assign out[488] = in[324];
    assign out[127] = in[325];
    assign out[40] = in[326];
    assign out[166] = in[327];
    assign out[275] = in[328];
    assign out[3] = in[329];
    assign out[312] = in[330];
    assign out[133] = in[331];
    assign out[110] = in[332];
    assign out[47] = in[333];
    assign out[148] = in[334];
    assign out[201] = in[335];
    assign out[175] = in[336];
    assign out[563] = in[337];
    assign out[577] = in[338];
    assign out[14] = in[339];
    assign out[289] = in[340];
    assign out[431] = in[341];
    assign out[632] = in[342];
    assign out[104] = in[343];
    assign out[122] = in[344];
    assign out[20] = in[345];
    assign out[433] = in[346];
    assign out[294] = in[347];
    assign out[189] = in[348];
    assign out[177] = in[349];
    assign out[297] = in[350];
    assign out[1] = in[351];
    assign out[530] = in[352];
    assign out[364] = in[353];
    assign out[206] = in[354];
    assign out[247] = in[355];
    assign out[94] = in[356];
    assign out[293] = in[357];
    assign out[210] = in[358];
    assign out[341] = in[359];
    assign out[278] = in[360];
    assign out[200] = in[361];
    assign out[398] = in[362];
    assign out[37] = in[363];
    assign out[390] = in[364];
    assign out[365] = in[365];
    assign out[379] = in[366];
    assign out[351] = in[367];
    assign out[495] = in[368];
    assign out[382] = in[369];
    assign out[145] = in[370];
    assign out[384] = in[371];
    assign out[250] = in[372];
    assign out[357] = in[373];
    assign out[138] = in[374];
    assign out[49] = in[375];
    assign out[554] = in[376];
    assign out[262] = in[377];
    assign out[540] = in[378];
    assign out[326] = in[379];
    assign out[82] = in[380];
    assign out[19] = in[381];
    assign out[331] = in[382];
    assign out[97] = in[383];
    assign out[514] = in[384];
    assign out[274] = in[385];
    assign out[529] = in[386];
    assign out[442] = in[387];
    assign out[277] = in[388];
    assign out[6] = in[389];
    assign out[533] = in[390];
    assign out[470] = in[391];
    assign out[302] = in[392];
    assign out[538] = in[393];
    assign out[368] = in[394];
    assign out[305] = in[395];
    assign out[438] = in[396];
    assign out[352] = in[397];
    assign out[626] = in[398];
    assign out[15] = in[399];
    assign out[320] = in[400];
    assign out[83] = in[401];
    assign out[457] = in[402];
    assign out[292] = in[403];
    assign out[22] = in[404];
    assign out[23] = in[405];
    assign out[136] = in[406];
    assign out[76] = in[407];
    assign out[617] = in[408];
    assign out[362] = in[409];
    assign out[272] = in[410];
    assign out[511] = in[411];
    assign out[606] = in[412];
    assign out[323] = in[413];
    assign out[183] = in[414];
    assign out[33] = in[415];
    assign out[354] = in[416];
    assign out[496] = in[417];
    assign out[373] = in[418];
    assign out[213] = in[419];
    assign out[520] = in[420];
    assign out[295] = in[421];
    assign out[525] = in[422];
    assign out[502] = in[423];
    assign out[396] = in[424];
    assign out[378] = in[425];
    assign out[61] = in[426];
    assign out[621] = in[427];
    assign out[366] = in[428];
    assign out[225] = in[429];
    assign out[445] = in[430];
    assign out[531] = in[431];
    assign out[57] = in[432];
    assign out[165] = in[433];
    assign out[534] = in[434];
    assign out[117] = in[435];
    assign out[261] = in[436];
    assign out[582] = in[437];
    assign out[592] = in[438];
    assign out[64] = in[439];
    assign out[58] = in[440];
    assign out[158] = in[441];
    assign out[221] = in[442];
    assign out[125] = in[443];
    assign out[149] = in[444];
    assign out[239] = in[445];
    assign out[215] = in[446];
    assign out[228] = in[447];
    assign out[548] = in[448];
    assign out[440] = in[449];
    assign out[428] = in[450];
    assign out[605] = in[451];
    assign out[535] = in[452];
    assign out[235] = in[453];
    assign out[59] = in[454];
    assign out[16] = in[455];
    assign out[539] = in[456];
    assign out[11] = in[457];
    assign out[314] = in[458];
    assign out[602] = in[459];
    assign out[451] = in[460];
    assign out[542] = in[461];
    assign out[67] = in[462];
    assign out[566] = in[463];
    assign out[194] = in[464];
    assign out[195] = in[465];
    assign out[355] = in[466];
    assign out[634] = in[467];
    assign out[198] = in[468];
    assign out[447] = in[469];
    assign out[461] = in[470];
    assign out[618] = in[471];
    assign out[444] = in[472];
    assign out[91] = in[473];
    assign out[638] = in[474];
    assign out[205] = in[475];
    assign out[111] = in[476];
    assign out[95] = in[477];
    assign out[578] = in[478];
    assign out[325] = in[479];
    assign out[458] = in[480];
    assign out[98] = in[481];
    assign out[612] = in[482];
    assign out[562] = in[483];
    assign out[100] = in[484];
    assign out[202] = in[485];
    assign out[552] = in[486];
    assign out[285] = in[487];
    assign out[633] = in[488];
    assign out[568] = in[489];
    assign out[468] = in[490];
    assign out[463] = in[491];
    assign out[381] = in[492];
    assign out[159] = in[493];
    assign out[472] = in[494];
    assign out[521] = in[495];
    assign out[147] = in[496];
    assign out[38] = in[497];
    assign out[259] = in[498];
    assign out[152] = in[499];
    assign out[603] = in[500];
    assign out[55] = in[501];
    assign out[517] = in[502];
    assign out[10] = in[503];
    assign out[482] = in[504];
    assign out[544] = in[505];
    assign out[484] = in[506];
    assign out[268] = in[507];
    assign out[126] = in[508];
    assign out[417] = in[509];
    assign out[501] = in[510];
    assign out[65] = in[511];
    assign out[121] = in[512];
    assign out[367] = in[513];
    assign out[230] = in[514];
    assign out[60] = in[515];
    assign out[422] = in[516];
    assign out[581] = in[517];
    assign out[151] = in[518];
    assign out[216] = in[519];
    assign out[340] = in[520];
    assign out[427] = in[521];
    assign out[174] = in[522];
    assign out[270] = in[523];
    assign out[412] = in[524];
    assign out[477] = in[525];
    assign out[105] = in[526];
    assign out[319] = in[527];
    assign out[629] = in[528];
    assign out[499] = in[529];
    assign out[436] = in[530];
    assign out[245] = in[531];
    assign out[241] = in[532];
    assign out[68] = in[533];
    assign out[504] = in[534];
    assign out[21] = in[535];
    assign out[86] = in[536];
    assign out[251] = in[537];
    assign out[137] = in[538];
    assign out[286] = in[539];
    assign out[190] = in[540];
    assign out[90] = in[541];
    assign out[430] = in[542];
    assign out[452] = in[543];
    assign out[337] = in[544];
    assign out[242] = in[545];
    assign out[196] = in[546];
    assign out[199] = in[547];
    assign out[500] = in[548];
    assign out[34] = in[549];
    assign out[279] = in[550];
    assign out[203] = in[551];
    assign out[616] = in[552];
    assign out[103] = in[553];
    assign out[39] = in[554];
    assign out[234] = in[555];
    assign out[508] = in[556];
    assign out[8] = in[557];
    assign out[510] = in[558];
    assign out[315] = in[559];
    assign out[407] = in[560];
    assign out[106] = in[561];
    assign out[13] = in[562];
    assign out[112] = in[563];
    assign out[35] = in[564];
    assign out[80] = in[565];
    assign out[115] = in[566];
    assign out[153] = in[567];
    assign out[413] = in[568];
    assign out[119] = in[569];
    assign out[78] = in[570];
    assign out[571] = in[571];
    assign out[478] = in[572];
    assign out[236] = in[573];
    assign out[595] = in[574];
    assign out[399] = in[575];
    assign out[400] = in[576];
    assign out[260] = in[577];
    assign out[599] = in[578];
    assign out[619] = in[579];
    assign out[88] = in[580];
    assign out[169] = in[581];
    assign out[311] = in[582];
    assign out[69] = in[583];
    assign out[92] = in[584];
    assign out[237] = in[585];
    assign out[231] = in[586];
    assign out[168] = in[587];
    assign out[139] = in[588];
    assign out[565] = in[589];
    assign out[75] = in[590];
    assign out[349] = in[591];
    assign out[107] = in[592];
    assign out[630] = in[593];
    assign out[102] = in[594];
    assign out[257] = in[595];
    assign out[507] = in[596];
    assign out[264] = in[597];
    assign out[486] = in[598];
    assign out[180] = in[599];
    assign out[469] = in[600];
    assign out[265] = in[601];
    assign out[171] = in[602];
    assign out[359] = in[603];
    assign out[476] = in[604];
    assign out[267] = in[605];
    assign out[298] = in[606];
    assign out[269] = in[607];
    assign out[416] = in[608];
    assign out[53] = in[609];
    assign out[586] = in[610];
    assign out[28] = in[611];
    assign out[306] = in[612];
    assign out[130] = in[613];
    assign out[590] = in[614];
    assign out[551] = in[615];
    assign out[281] = in[616];
    assign out[309] = in[617];
    assign out[99] = in[618];
    assign out[402] = in[619];
    assign out[303] = in[620];
    assign out[350] = in[621];
    assign out[515] = in[622];
    assign out[288] = in[623];
    assign out[141] = in[624];
    assign out[372] = in[625];
    assign out[386] = in[626];
    assign out[208] = in[627];
    assign out[473] = in[628];
    assign out[51] = in[629];
    assign out[258] = in[630];
    assign out[182] = in[631];
    assign out[324] = in[632];
    assign out[248] = in[633];
    assign out[610] = in[634];
    assign out[611] = in[635];
    assign out[460] = in[636];
    assign out[118] = in[637];
    assign out[421] = in[638];
    assign out[301] = in[639];
endmodule

module encrypt_4rotation_helper(in, out);
    input [63:0] in;
    output [63:0] out;
    assign out = {in[58:0], in[63:59]} ^ {in[53:0], in[63:54]} ^ {in[5:0], in[63:6]} ^ {in[30:0], in[63:31]} ^ {in[2:0], in[63:3]} ^ {in[59:0], in[63:60]};
endmodule

module encrypt_4apply_rotations(in, out);
    input [639:0] in;
    output [639:0] out;
    wire [639:0] rot;
    encrypt_4rotation_helper rot0inst(in[63:0], rot[63:0]);
    encrypt_4rotation_helper rot1inst(in[127:64], rot[127:64]);
    encrypt_4rotation_helper rot2inst(in[191:128], rot[191:128]);
    encrypt_4rotation_helper rot3inst(in[255:192], rot[255:192]);
    encrypt_4rotation_helper rot4inst(in[319:256], rot[319:256]);
    encrypt_4rotation_helper rot5inst(in[383:320], rot[383:320]);
    encrypt_4rotation_helper rot6inst(in[447:384], rot[447:384]);
    encrypt_4rotation_helper rot7inst(in[511:448], rot[511:448]);
    encrypt_4rotation_helper rot8inst(in[575:512], rot[575:512]);
    encrypt_4rotation_helper rot9inst(in[639:576], rot[639:576]);
    assign out = rot ^ {in[63:0], in[639:64]};
endmodule

module encrypt_4apply_round_key(key, in, out);
    input [9:0] key;
    input [639:0] in;
    output [639:0] out;
    assign out[0] = in[0] ^ key[0];
    assign out[63:1] = in[63:1];
    assign out[64] = in[64] ^ key[1];
    assign out[127:65] = in[127:65];
    assign out[128] = in[128] ^ key[2];
    assign out[191:129] = in[191:129];
    assign out[192] = in[192] ^ key[3];
    assign out[255:193] = in[255:193];
    assign out[256] = in[256] ^ key[4];
    assign out[319:257] = in[319:257];
    assign out[320] = in[320] ^ key[5];
    assign out[383:321] = in[383:321];
    assign out[384] = in[384] ^ key[6];
    assign out[447:385] = in[447:385];
    assign out[448] = in[448] ^ key[7];
    assign out[511:449] = in[511:449];
    assign out[512] = in[512] ^ key[8];
    assign out[575:513] = in[575:513];
    assign out[576] = in[576] ^ key[9];
    assign out[639:577] = in[639:577];
endmodule

module encrypt_4full_round(clk, roundkey, in, out);
    input clk;
    input [9:0] roundkey;
    input [639:0] in;
    output [639:0] out;
    wire [639:0] mid[0:3];
    encrypt_4apply_pbox0 pbox0inst(in, mid[0]);
    encrypt_4apply_sboxes sboxes(clk, mid[0], mid[1]);
    encrypt_4apply_pbox1 pbox1inst(mid[1], mid[2]);
    encrypt_4apply_rotations rotations(mid[2], mid[3]);
    encrypt_4apply_round_key keys(roundkey, mid[3], out);
endmodule

module encrypt_4get_round_key0(clk, period, key);
    input clk;
    input [1:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        2'h0: key <= 10'h3e9;
        2'h1: key <= 10'h394;
        2'h2: key <= 10'h3f0;
        2'h3: key <= 10'h104;
    endcase
    end
endmodule

module encrypt_4get_round_key1(clk, period, key);
    input clk;
    input [1:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        2'h0: key <= 10'h201;
        2'h1: key <= 10'h0da;
        2'h2: key <= 10'h36d;
        2'h3: key <= 10'h178;
    endcase
    end
endmodule

module encrypt_4get_round_key2(clk, period, key);
    input clk;
    input [1:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        2'h0: key <= 10'h097;
        2'h1: key <= 10'h0d7;
        2'h2: key <= 10'h35c;
        2'h3: key <= 10'h0aa;
    endcase
    end
endmodule

module encrypt_4get_round_key3(clk, period, key);
    input clk;
    input [1:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        2'h0: key <= 10'h116;
        2'h1: key <= 10'h321;
        2'h2: key <= 10'h14f;
        2'h3: key <= 10'h20a;
    endcase
    end
endmodule

module encrypt_4get_round_key4(clk, period, key);
    input clk;
    input [1:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        2'h0: key <= 10'h131;
        2'h1: key <= 10'h123;
        2'h2: key <= 10'h1dd;
        2'h3: key <= 10'h1bf;
    endcase
    end
endmodule

module encrypt_4get_round_key5(clk, period, key);
    input clk;
    input [1:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        2'h0: key <= 10'h353;
        2'h1: key <= 10'h151;
        2'h2: key <= 10'h14c;
        2'h3: key <= 10'h2ac;
    endcase
    end
endmodule

module encrypt_4get_round_key6(clk, period, key);
    input clk;
    input [1:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        2'h0: key <= 10'h010;
        2'h1: key <= 10'h3ae;
        2'h2: key <= 10'h2fa;
        2'h3: key <= 10'h2d9;
    endcase
    end
endmodule

module encrypt_4get_round_key7(clk, period, key);
    input clk;
    input [1:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        2'h0: key <= 10'h046;
        2'h1: key <= 10'h354;
        2'h2: key <= 10'h249;
        2'h3: key <= 10'h31c;
    endcase
    end
endmodule

module encrypt_4get_round_key8(clk, period, key);
    input clk;
    input [1:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        2'h0: key <= 10'h3ee;
        2'h1: key <= 10'h2c6;
        2'h2: key <= 10'h14b;
        2'h3: key <= 10'h293;
    endcase
    end
endmodule

module encrypt_4get_round_key9(clk, period, key);
    input clk;
    input [1:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        2'h0: key <= 10'h042;
        2'h1: key <= 10'h3ba;
        2'h2: key <= 10'h304;
        2'h3: key <= 10'h206;
    endcase
    end
endmodule

module encrypt_4get_round_key10(clk, period, key);
    input clk;
    input [1:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        2'h0: key <= 10'h004;
        2'h1: key <= 10'h239;
        2'h2: key <= 10'h1c1;
        2'h3: key <= 10'h2b9;
    endcase
    end
endmodule

module encrypt_4get_round_key11(clk, period, key);
    input clk;
    input [1:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        2'h0: key <= 10'h069;
        2'h1: key <= 10'h0d6;
        2'h2: key <= 10'h2e4;
        2'h3: key <= 10'h170;
    endcase
    end
endmodule

module encrypt_4get_round_key12(clk, period, key);
    input clk;
    input [1:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        2'h0: key <= 10'h06e;
        2'h1: key <= 10'h29a;
        2'h2: key <= 10'h35c;
        2'h3: key <= 10'h31f;
    endcase
    end
endmodule

module encrypt_4get_round_key13(clk, period, key);
    input clk;
    input [1:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        2'h0: key <= 10'h239;
        2'h1: key <= 10'h288;
        2'h2: key <= 10'h251;
        2'h3: key <= 10'h36c;
    endcase
    end
endmodule

module encrypt_4get_round_key14(clk, period, key);
    input clk;
    input [1:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        2'h0: key <= 10'h1aa;
        2'h1: key <= 10'h242;
        2'h2: key <= 10'h317;
        2'h3: key <= 10'h23b;
    endcase
    end
endmodule

module encrypt_4get_round_key15(clk, period, key);
    input clk;
    input [1:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        2'h0: key <= 10'h1ff;
        2'h1: key <= 10'h348;
        2'h2: key <= 10'h11e;
        2'h3: key <= 10'h186;
    endcase
    end
endmodule

module encrypt_4get_round_key16(clk, period, key);
    input clk;
    input [1:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        2'h0: key <= 10'h0b6;
        2'h1: key <= 10'h2be;
        2'h2: key <= 10'h250;
        2'h3: key <= 10'h3c9;
    endcase
    end
endmodule

module encrypt_4get_round_key17(clk, period, key);
    input clk;
    input [1:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        2'h0: key <= 10'h368;
        2'h1: key <= 10'h171;
        2'h2: key <= 10'h2dc;
        2'h3: key <= 10'h161;
    endcase
    end
endmodule

module encrypt_4get_round_key18(clk, period, key);
    input clk;
    input [1:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        2'h0: key <= 10'h127;
        2'h1: key <= 10'h159;
        2'h2: key <= 10'h1fd;
        2'h3: key <= 10'h006;
    endcase
    end
endmodule

module encrypt_4get_round_key19(clk, period, key);
    input clk;
    input [1:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        2'h0: key <= 10'h1b3;
        2'h1: key <= 10'h390;
        2'h2: key <= 10'h185;
        2'h3: key <= 10'h1d5;
    endcase
    end
endmodule

module encrypt_4get_round_key20(clk, period, key);
    input clk;
    input [1:0] period;
    output [9:0] key;
    reg [9:0] key;
    always @(posedge clk) begin
    case (period)
        2'h0: key <= 10'h314;
        2'h1: key <= 10'h103;
        2'h2: key <= 10'h1e7;
        2'h3: key <= 10'h0bb;
    endcase
    end
endmodule

module encrypt_4encrypt_loop(clk, in, read, out, write);
    input clk;
    input [639:0] in;
    input read;
    output reg [639:0] out;
    output write;
    reg [639:0] state[21:0];
    wire [639:0] next[21:0];
    always @(posedge clk) state[1] <= next[0];
    always @(posedge clk) state[2] <= next[1];
    always @(posedge clk) state[3] <= next[2];
    always @(posedge clk) state[4] <= next[3];
    always @(posedge clk) state[5] <= next[4];
    always @(posedge clk) state[6] <= next[5];
    always @(posedge clk) state[7] <= next[6];
    always @(posedge clk) state[8] <= next[7];
    always @(posedge clk) state[9] <= next[8];
    always @(posedge clk) state[10] <= next[9];
    always @(posedge clk) state[11] <= next[10];
    always @(posedge clk) state[12] <= next[11];
    always @(posedge clk) state[13] <= next[12];
    always @(posedge clk) state[14] <= next[13];
    always @(posedge clk) state[15] <= next[14];
    always @(posedge clk) state[16] <= next[15];
    always @(posedge clk) state[17] <= next[16];
    always @(posedge clk) state[18] <= next[17];
    always @(posedge clk) state[19] <= next[18];
    always @(posedge clk) state[20] <= next[19];
    always @(posedge clk) state[21] <= next[20];
    assign next[21] = state[21];
    wire [9:0] roundkey[20:0];
    reg [1:0] period[42:0];
    always @(posedge clk) period[1] <= period[0];
    always @(posedge clk) period[2] <= period[1];
    always @(posedge clk) period[3] <= period[2];
    always @(posedge clk) period[4] <= period[3];
    always @(posedge clk) period[5] <= period[4];
    always @(posedge clk) period[6] <= period[5];
    always @(posedge clk) period[7] <= period[6];
    always @(posedge clk) period[8] <= period[7];
    always @(posedge clk) period[9] <= period[8];
    always @(posedge clk) period[10] <= period[9];
    always @(posedge clk) period[11] <= period[10];
    always @(posedge clk) period[12] <= period[11];
    always @(posedge clk) period[13] <= period[12];
    always @(posedge clk) period[14] <= period[13];
    always @(posedge clk) period[15] <= period[14];
    always @(posedge clk) period[16] <= period[15];
    always @(posedge clk) period[17] <= period[16];
    always @(posedge clk) period[18] <= period[17];
    always @(posedge clk) period[19] <= period[18];
    always @(posedge clk) period[20] <= period[19];
    always @(posedge clk) period[21] <= period[20];
    always @(posedge clk) period[22] <= period[21];
    always @(posedge clk) period[23] <= period[22];
    always @(posedge clk) period[24] <= period[23];
    always @(posedge clk) period[25] <= period[24];
    always @(posedge clk) period[26] <= period[25];
    always @(posedge clk) period[27] <= period[26];
    always @(posedge clk) period[28] <= period[27];
    always @(posedge clk) period[29] <= period[28];
    always @(posedge clk) period[30] <= period[29];
    always @(posedge clk) period[31] <= period[30];
    always @(posedge clk) period[32] <= period[31];
    always @(posedge clk) period[33] <= period[32];
    always @(posedge clk) period[34] <= period[33];
    always @(posedge clk) period[35] <= period[34];
    always @(posedge clk) period[36] <= period[35];
    always @(posedge clk) period[37] <= period[36];
    always @(posedge clk) period[38] <= period[37];
    always @(posedge clk) period[39] <= period[38];
    always @(posedge clk) period[40] <= period[39];
    always @(posedge clk) period[41] <= period[40];
    always @(posedge clk) period[42] <= period[41];
    encrypt_4get_round_key0 get_key0(clk, period[0], roundkey[0]);
    encrypt_4full_round round0(clk, roundkey[0], state[0], next[0]);
    encrypt_4get_round_key1 get_key1(clk, period[2], roundkey[1]);
    encrypt_4full_round round1(clk, roundkey[1], state[1], next[1]);
    encrypt_4get_round_key2 get_key2(clk, period[4], roundkey[2]);
    encrypt_4full_round round2(clk, roundkey[2], state[2], next[2]);
    encrypt_4get_round_key3 get_key3(clk, period[6], roundkey[3]);
    encrypt_4full_round round3(clk, roundkey[3], state[3], next[3]);
    encrypt_4get_round_key4 get_key4(clk, period[8], roundkey[4]);
    encrypt_4full_round round4(clk, roundkey[4], state[4], next[4]);
    encrypt_4get_round_key5 get_key5(clk, period[10], roundkey[5]);
    encrypt_4full_round round5(clk, roundkey[5], state[5], next[5]);
    encrypt_4get_round_key6 get_key6(clk, period[12], roundkey[6]);
    encrypt_4full_round round6(clk, roundkey[6], state[6], next[6]);
    encrypt_4get_round_key7 get_key7(clk, period[14], roundkey[7]);
    encrypt_4full_round round7(clk, roundkey[7], state[7], next[7]);
    encrypt_4get_round_key8 get_key8(clk, period[16], roundkey[8]);
    encrypt_4full_round round8(clk, roundkey[8], state[8], next[8]);
    encrypt_4get_round_key9 get_key9(clk, period[18], roundkey[9]);
    encrypt_4full_round round9(clk, roundkey[9], state[9], next[9]);
    encrypt_4get_round_key10 get_key10(clk, period[20], roundkey[10]);
    encrypt_4full_round round10(clk, roundkey[10], state[10], next[10]);
    encrypt_4get_round_key11 get_key11(clk, period[22], roundkey[11]);
    encrypt_4full_round round11(clk, roundkey[11], state[11], next[11]);
    encrypt_4get_round_key12 get_key12(clk, period[24], roundkey[12]);
    encrypt_4full_round round12(clk, roundkey[12], state[12], next[12]);
    encrypt_4get_round_key13 get_key13(clk, period[26], roundkey[13]);
    encrypt_4full_round round13(clk, roundkey[13], state[13], next[13]);
    encrypt_4get_round_key14 get_key14(clk, period[28], roundkey[14]);
    encrypt_4full_round round14(clk, roundkey[14], state[14], next[14]);
    encrypt_4get_round_key15 get_key15(clk, period[30], roundkey[15]);
    encrypt_4full_round round15(clk, roundkey[15], state[15], next[15]);
    encrypt_4get_round_key16 get_key16(clk, period[32], roundkey[16]);
    encrypt_4full_round round16(clk, roundkey[16], state[16], next[16]);
    encrypt_4get_round_key17 get_key17(clk, period[34], roundkey[17]);
    encrypt_4full_round round17(clk, roundkey[17], state[17], next[17]);
    encrypt_4get_round_key18 get_key18(clk, period[36], roundkey[18]);
    encrypt_4full_round round18(clk, roundkey[18], state[18], next[18]);
    encrypt_4get_round_key19 get_key19(clk, period[38], roundkey[19]);
    encrypt_4full_round round19(clk, roundkey[19], state[19], next[19]);
    encrypt_4get_round_key20 get_key20(clk, period[40], roundkey[20]);
    encrypt_4full_round round20(clk, roundkey[20], state[20], next[20]);
    always @(posedge clk) begin
        if (read)
        begin
            period[0] <= 0;
            state[0] <= in;
        end
        else
        begin
            period[0] <= period[42]+1;
            state[0] <= next[21];
        end
        out <= next[20];
    end
    reg [171:0] progress;
    initial progress = 172'h0;
    always @(posedge clk) progress[0] <= read;
    always @(posedge clk) progress[1] <= progress[0];
    always @(posedge clk) progress[2] <= progress[1];
    always @(posedge clk) progress[3] <= progress[2];
    always @(posedge clk) progress[4] <= progress[3];
    always @(posedge clk) progress[5] <= progress[4];
    always @(posedge clk) progress[6] <= progress[5];
    always @(posedge clk) progress[7] <= progress[6];
    always @(posedge clk) progress[8] <= progress[7];
    always @(posedge clk) progress[9] <= progress[8];
    always @(posedge clk) progress[10] <= progress[9];
    always @(posedge clk) progress[11] <= progress[10];
    always @(posedge clk) progress[12] <= progress[11];
    always @(posedge clk) progress[13] <= progress[12];
    always @(posedge clk) progress[14] <= progress[13];
    always @(posedge clk) progress[15] <= progress[14];
    always @(posedge clk) progress[16] <= progress[15];
    always @(posedge clk) progress[17] <= progress[16];
    always @(posedge clk) progress[18] <= progress[17];
    always @(posedge clk) progress[19] <= progress[18];
    always @(posedge clk) progress[20] <= progress[19];
    always @(posedge clk) progress[21] <= progress[20];
    always @(posedge clk) progress[22] <= progress[21];
    always @(posedge clk) progress[23] <= progress[22];
    always @(posedge clk) progress[24] <= progress[23];
    always @(posedge clk) progress[25] <= progress[24];
    always @(posedge clk) progress[26] <= progress[25];
    always @(posedge clk) progress[27] <= progress[26];
    always @(posedge clk) progress[28] <= progress[27];
    always @(posedge clk) progress[29] <= progress[28];
    always @(posedge clk) progress[30] <= progress[29];
    always @(posedge clk) progress[31] <= progress[30];
    always @(posedge clk) progress[32] <= progress[31];
    always @(posedge clk) progress[33] <= progress[32];
    always @(posedge clk) progress[34] <= progress[33];
    always @(posedge clk) progress[35] <= progress[34];
    always @(posedge clk) progress[36] <= progress[35];
    always @(posedge clk) progress[37] <= progress[36];
    always @(posedge clk) progress[38] <= progress[37];
    always @(posedge clk) progress[39] <= progress[38];
    always @(posedge clk) progress[40] <= progress[39];
    always @(posedge clk) progress[41] <= progress[40];
    always @(posedge clk) progress[42] <= progress[41];
    always @(posedge clk) progress[43] <= progress[42];
    always @(posedge clk) progress[44] <= progress[43];
    always @(posedge clk) progress[45] <= progress[44];
    always @(posedge clk) progress[46] <= progress[45];
    always @(posedge clk) progress[47] <= progress[46];
    always @(posedge clk) progress[48] <= progress[47];
    always @(posedge clk) progress[49] <= progress[48];
    always @(posedge clk) progress[50] <= progress[49];
    always @(posedge clk) progress[51] <= progress[50];
    always @(posedge clk) progress[52] <= progress[51];
    always @(posedge clk) progress[53] <= progress[52];
    always @(posedge clk) progress[54] <= progress[53];
    always @(posedge clk) progress[55] <= progress[54];
    always @(posedge clk) progress[56] <= progress[55];
    always @(posedge clk) progress[57] <= progress[56];
    always @(posedge clk) progress[58] <= progress[57];
    always @(posedge clk) progress[59] <= progress[58];
    always @(posedge clk) progress[60] <= progress[59];
    always @(posedge clk) progress[61] <= progress[60];
    always @(posedge clk) progress[62] <= progress[61];
    always @(posedge clk) progress[63] <= progress[62];
    always @(posedge clk) progress[64] <= progress[63];
    always @(posedge clk) progress[65] <= progress[64];
    always @(posedge clk) progress[66] <= progress[65];
    always @(posedge clk) progress[67] <= progress[66];
    always @(posedge clk) progress[68] <= progress[67];
    always @(posedge clk) progress[69] <= progress[68];
    always @(posedge clk) progress[70] <= progress[69];
    always @(posedge clk) progress[71] <= progress[70];
    always @(posedge clk) progress[72] <= progress[71];
    always @(posedge clk) progress[73] <= progress[72];
    always @(posedge clk) progress[74] <= progress[73];
    always @(posedge clk) progress[75] <= progress[74];
    always @(posedge clk) progress[76] <= progress[75];
    always @(posedge clk) progress[77] <= progress[76];
    always @(posedge clk) progress[78] <= progress[77];
    always @(posedge clk) progress[79] <= progress[78];
    always @(posedge clk) progress[80] <= progress[79];
    always @(posedge clk) progress[81] <= progress[80];
    always @(posedge clk) progress[82] <= progress[81];
    always @(posedge clk) progress[83] <= progress[82];
    always @(posedge clk) progress[84] <= progress[83];
    always @(posedge clk) progress[85] <= progress[84];
    always @(posedge clk) progress[86] <= progress[85];
    always @(posedge clk) progress[87] <= progress[86];
    always @(posedge clk) progress[88] <= progress[87];
    always @(posedge clk) progress[89] <= progress[88];
    always @(posedge clk) progress[90] <= progress[89];
    always @(posedge clk) progress[91] <= progress[90];
    always @(posedge clk) progress[92] <= progress[91];
    always @(posedge clk) progress[93] <= progress[92];
    always @(posedge clk) progress[94] <= progress[93];
    always @(posedge clk) progress[95] <= progress[94];
    always @(posedge clk) progress[96] <= progress[95];
    always @(posedge clk) progress[97] <= progress[96];
    always @(posedge clk) progress[98] <= progress[97];
    always @(posedge clk) progress[99] <= progress[98];
    always @(posedge clk) progress[100] <= progress[99];
    always @(posedge clk) progress[101] <= progress[100];
    always @(posedge clk) progress[102] <= progress[101];
    always @(posedge clk) progress[103] <= progress[102];
    always @(posedge clk) progress[104] <= progress[103];
    always @(posedge clk) progress[105] <= progress[104];
    always @(posedge clk) progress[106] <= progress[105];
    always @(posedge clk) progress[107] <= progress[106];
    always @(posedge clk) progress[108] <= progress[107];
    always @(posedge clk) progress[109] <= progress[108];
    always @(posedge clk) progress[110] <= progress[109];
    always @(posedge clk) progress[111] <= progress[110];
    always @(posedge clk) progress[112] <= progress[111];
    always @(posedge clk) progress[113] <= progress[112];
    always @(posedge clk) progress[114] <= progress[113];
    always @(posedge clk) progress[115] <= progress[114];
    always @(posedge clk) progress[116] <= progress[115];
    always @(posedge clk) progress[117] <= progress[116];
    always @(posedge clk) progress[118] <= progress[117];
    always @(posedge clk) progress[119] <= progress[118];
    always @(posedge clk) progress[120] <= progress[119];
    always @(posedge clk) progress[121] <= progress[120];
    always @(posedge clk) progress[122] <= progress[121];
    always @(posedge clk) progress[123] <= progress[122];
    always @(posedge clk) progress[124] <= progress[123];
    always @(posedge clk) progress[125] <= progress[124];
    always @(posedge clk) progress[126] <= progress[125];
    always @(posedge clk) progress[127] <= progress[126];
    always @(posedge clk) progress[128] <= progress[127];
    always @(posedge clk) progress[129] <= progress[128];
    always @(posedge clk) progress[130] <= progress[129];
    always @(posedge clk) progress[131] <= progress[130];
    always @(posedge clk) progress[132] <= progress[131];
    always @(posedge clk) progress[133] <= progress[132];
    always @(posedge clk) progress[134] <= progress[133];
    always @(posedge clk) progress[135] <= progress[134];
    always @(posedge clk) progress[136] <= progress[135];
    always @(posedge clk) progress[137] <= progress[136];
    always @(posedge clk) progress[138] <= progress[137];
    always @(posedge clk) progress[139] <= progress[138];
    always @(posedge clk) progress[140] <= progress[139];
    always @(posedge clk) progress[141] <= progress[140];
    always @(posedge clk) progress[142] <= progress[141];
    always @(posedge clk) progress[143] <= progress[142];
    always @(posedge clk) progress[144] <= progress[143];
    always @(posedge clk) progress[145] <= progress[144];
    always @(posedge clk) progress[146] <= progress[145];
    always @(posedge clk) progress[147] <= progress[146];
    always @(posedge clk) progress[148] <= progress[147];
    always @(posedge clk) progress[149] <= progress[148];
    always @(posedge clk) progress[150] <= progress[149];
    always @(posedge clk) progress[151] <= progress[150];
    always @(posedge clk) progress[152] <= progress[151];
    always @(posedge clk) progress[153] <= progress[152];
    always @(posedge clk) progress[154] <= progress[153];
    always @(posedge clk) progress[155] <= progress[154];
    always @(posedge clk) progress[156] <= progress[155];
    always @(posedge clk) progress[157] <= progress[156];
    always @(posedge clk) progress[158] <= progress[157];
    always @(posedge clk) progress[159] <= progress[158];
    always @(posedge clk) progress[160] <= progress[159];
    always @(posedge clk) progress[161] <= progress[160];
    always @(posedge clk) progress[162] <= progress[161];
    always @(posedge clk) progress[163] <= progress[162];
    always @(posedge clk) progress[164] <= progress[163];
    always @(posedge clk) progress[165] <= progress[164];
    always @(posedge clk) progress[166] <= progress[165];
    always @(posedge clk) progress[167] <= progress[166];
    always @(posedge clk) progress[168] <= progress[167];
    always @(posedge clk) progress[169] <= progress[168];
    always @(posedge clk) progress[170] <= progress[169];
    always @(posedge clk) progress[171] <= progress[170];
    assign write = progress[171];
endmodule

module encrypt_4encrypt(clk, in, read, out, write);
    localparam THROUGHPUT = 4;
    input clk;
    input [639:0] in;
    input read;
    output [639:0] out;
    output write;
    reg [1:0] progress;
    initial progress = 2'h0;
    reg [639:0] state[1:0];
    wire [639:0] next;
    encrypt_4pre_mix premixer(state[0], next);
    encrypt_4encrypt_loop crypter(clk, state[1], progress[1], out, write);
    always @(posedge clk) begin
        progress[0] <= read;
        progress[1] <= progress[0];
        state[0] <= in;
        state[1] <= next;
    end
endmodule
